.include TSMC_180nm.txt
.param SUPPLY=1.8
.param LAMBDA=0.09u
.param w = {20*LAMBDA}
.param width_P={2*w}
.param width_N={2*w}
.param width_P_i = (LAMBDA*50)
.param width_N_i = (LAMBDA*20)
.global gnd vdd

Vdd	vdd	gnd	'SUPPLY'

vin1 A0 0 pulse 0 1.8 0n 100p 100p 19.9n 40n
vin2 A1 0 pulse 0 1.8 0n 100p 100p 19.9n 40n
vin3 A2 0 pulse 0 1.8 0n 100p 100p 19.9n 40n
vin4 A3 0 pulse 0 1.8 0n 100p 100p 19.9n 40n

vin5 B0 0 pulse 0 1.8 0n 100p 100p 49.9n 100n
vin6 B1 0 pulse 0 1.8 0n 100p 100p 49.9n 100n
vin7 B2 0 pulse 0 1.8 0n 100p 100p 49.9n 100n
vin8 B3 0 pulse 0 1.8 0n 100p 100p 49.9n 100n



.subckt nand A B out vdd gnd
M1      out       A       k     gnd  CMOSN   W={width_N}   L={2*LAMBDA}
+ AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N} AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}

M2      out       A       vdd     vdd  CMOSP   W={width_P}   L={2*LAMBDA}
+ AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P} AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}

M3      k       B       gnd     gnd  CMOSN   W={width_N}   L={2*LAMBDA}
+ AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N} AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}

M4      out       B       vdd     vdd  CMOSP   W={width_P}   L={2*LAMBDA}
+ AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P} AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}
.ends nand

.subckt inv yi xi vdd gnd
M1      yi       xi       gnd     gnd  CMOSN   W={width_N_i}   L={2*LAMBDA}
+ AS={5*width_N_i*LAMBDA} PS={10*LAMBDA+2*width_N_i} AD={5*width_N_i*LAMBDA} PD={10*LAMBDA+2*width_N}
M2      yi       xi       vdd     vdd  CMOSP   W={width_P_i}   L={2*LAMBDA}
+ AS={5*width_P_i*LAMBDA} PS={10*LAMBDA+2*width_P_i} AD={5*width_P_i*LAMBDA} PD={10*LAMBDA+2*width_P_i}
.ends inv


***********XOR gate*******************
.subckt xor dma dmb outx vdd gnd
xx1 dma dmb outx1 vdd gnd nand
xx2 dma outx1 outx2 vdd gnd nand
xx3 dmb outx1 outx3 vdd gnd nand
xx4 outx2 outx3 outx vdd gnd nand
.ends xor  

**************AND GATE*******************
.subckt and_g in1 in2 aout vdd gnd
xx5 in1 in2 out_nan vdd gnd nand
xx6 aout out_nan  vdd gnd inv
.ends and_g

*****************OR GATE*****************
.subckt or_g inn1 inn2 orout vdd gnd
xx7 ou1 inn1 vdd gnd inv
xx8 ou2 inn2 vdd gnd inv
xx9 ou1 ou2 orout vdd gnd nand
.ends or_g


**********************Generate*********************

x140 A0 B0   g0 vdd gnd and_g
x141 A1 B1  g1 vdd gnd and_g
x142 A2 B2  g2 vdd gnd and_g
x143 A3 B3  g3 vdd gnd and_g

**********************Propagate********************
x144 A0   B0   p0 vdd gnd xor
x145 A1  B1  p1 vdd gnd xor
x146 A2  B2  p2 vdd gnd xor
x147 A3  B3  p3 vdd gnd xor



.tran 0.1n 200n

.control
set hcopypscolor = 1
set color0=white
set color1=black

run
set curplottitle="Ayush-2020122001"

*plot v(s_bar)
*plot v(clk)
plot v(A0) v(B0)
plot v(p0)
plot v(g0)
set hcopypscolor = 1
hardcopy propagate.eps v(p0)
hardcopy input.eps v(A0) v(B0)
hardcopy generate.eps v(g0)
.endc
