magic
tech scmos
timestamp 1619456195
<< nwell >>
rect 15 4173 71 4270
rect 265 4173 321 4270
rect 345 4173 401 4270
rect 595 4173 651 4270
rect 258 4118 337 4143
rect 266 3997 322 4094
rect 266 3871 322 3968
rect 346 3871 402 3968
rect 2222 3864 2319 3920
rect 1170 3610 1249 3635
rect 2222 3614 2319 3670
rect 2524 3615 2621 3671
rect 1178 3479 1234 3576
rect 2222 3534 2319 3590
rect 2349 3527 2374 3606
rect 2398 3535 2495 3591
rect 2524 3535 2621 3591
rect 1170 3436 1249 3461
rect 1923 3449 2020 3505
rect 1178 3314 1234 3411
rect 1799 3370 1896 3426
rect 1923 3369 2020 3425
rect 2038 3369 2135 3425
rect 15 3216 71 3313
rect 265 3216 321 3313
rect 345 3216 401 3313
rect 595 3216 651 3313
rect 1171 3277 1250 3302
rect 2222 3284 2319 3340
rect 2222 3204 2319 3260
rect 258 3161 337 3186
rect 266 3040 322 3137
rect 729 3091 826 3147
rect 853 3092 950 3148
rect 968 3092 1065 3148
rect 1187 3093 1243 3190
rect 853 3012 950 3068
rect 1180 3056 1259 3081
rect 266 2914 322 3011
rect 346 2914 402 3011
rect 15 2737 71 2834
rect 265 2737 321 2834
rect 345 2737 401 2834
rect 595 2737 651 2834
rect 714 2798 770 2895
rect 1188 2888 1244 2985
rect 1799 2971 1896 3027
rect 1923 2972 2020 3028
rect 2038 2972 2135 3028
rect 2222 2954 2319 3010
rect 2524 2955 2621 3011
rect 1923 2892 2020 2948
rect 1181 2851 1260 2876
rect 2222 2874 2319 2930
rect 2349 2867 2374 2946
rect 2398 2875 2495 2931
rect 2524 2875 2621 2931
rect 698 2761 777 2786
rect 1181 2770 1260 2795
rect 258 2682 337 2707
rect 266 2561 322 2658
rect 698 2631 777 2656
rect 1189 2639 1245 2736
rect 1298 2720 1377 2745
rect 266 2435 322 2532
rect 346 2435 402 2532
rect 714 2522 770 2619
rect 1181 2596 1260 2621
rect 1313 2589 1369 2686
rect 2222 2624 2319 2680
rect 1298 2546 1377 2571
rect 2222 2544 2319 2600
rect 15 2258 71 2355
rect 265 2258 321 2355
rect 345 2258 401 2355
rect 595 2258 651 2355
rect 853 2349 950 2405
rect 1361 2365 1440 2390
rect 729 2270 826 2326
rect 853 2269 950 2325
rect 968 2269 1065 2325
rect 1083 2269 1180 2325
rect 1192 2262 1217 2341
rect 1376 2234 1432 2331
rect 1923 2323 2020 2379
rect 1799 2244 1896 2300
rect 1923 2243 2020 2299
rect 2038 2243 2135 2299
rect 2222 2294 2319 2350
rect 2524 2295 2621 2351
rect 258 2203 337 2228
rect 1361 2191 1440 2216
rect 1632 2195 1711 2220
rect 2222 2214 2319 2270
rect 2349 2207 2374 2286
rect 2398 2215 2495 2271
rect 2524 2215 2621 2271
rect 266 2082 322 2179
rect 1365 2130 1444 2155
rect 266 1956 322 2053
rect 346 1956 402 2053
rect 729 1965 826 2021
rect 853 1966 950 2022
rect 968 1966 1065 2022
rect 1083 2019 1180 2075
rect 1192 2003 1217 2082
rect 1380 1999 1436 2096
rect 1640 2064 1696 2161
rect 1632 2021 1711 2046
rect 853 1886 950 1942
rect 1083 1923 1180 1979
rect 1192 1916 1217 1995
rect 1365 1956 1444 1981
rect 2222 1964 2319 2020
rect 15 1779 71 1876
rect 265 1779 321 1876
rect 345 1779 401 1876
rect 595 1779 651 1876
rect 1799 1845 1896 1901
rect 1923 1846 2020 1902
rect 2038 1846 2135 1902
rect 2222 1884 2319 1940
rect 258 1724 337 1749
rect 266 1603 322 1700
rect 714 1672 770 1769
rect 1923 1766 2020 1822
rect 698 1635 777 1660
rect 1080 1636 1177 1692
rect 1189 1620 1214 1699
rect 2222 1634 2319 1690
rect 2524 1635 2621 1691
rect 1458 1594 1537 1619
rect 266 1477 322 1574
rect 346 1477 402 1574
rect 1076 1435 1173 1491
rect 1185 1419 1210 1498
rect 1473 1463 1529 1560
rect 2222 1554 2319 1610
rect 2349 1547 2374 1626
rect 2398 1555 2495 1611
rect 2524 1555 2621 1611
rect 1458 1420 1537 1445
rect 1729 1424 1808 1449
rect 15 1300 71 1397
rect 265 1300 321 1397
rect 345 1300 401 1397
rect 595 1300 651 1397
rect 1076 1341 1173 1397
rect 1185 1334 1210 1413
rect 1462 1359 1541 1384
rect 258 1245 337 1270
rect 1477 1228 1533 1325
rect 1737 1293 1793 1390
rect 2222 1304 2319 1360
rect 1729 1250 1808 1275
rect 2222 1224 2319 1280
rect 266 1124 322 1221
rect 1462 1185 1541 1210
rect 1720 1162 1799 1187
rect 266 998 322 1095
rect 346 998 402 1095
rect 1076 1062 1173 1118
rect 1185 1046 1210 1125
rect 1728 1031 1784 1128
rect 1720 988 1799 1013
rect 2222 974 2319 1030
rect 2524 975 2621 1031
rect 15 821 71 918
rect 265 821 321 918
rect 345 821 401 918
rect 595 821 651 918
rect 2222 894 2319 950
rect 2349 887 2374 966
rect 2398 895 2495 951
rect 2524 895 2621 951
rect 258 766 337 791
rect 266 645 322 742
rect 2222 644 2319 700
rect 266 519 322 616
rect 346 519 402 616
rect 15 342 71 439
rect 265 342 321 439
rect 345 342 401 439
rect 595 342 651 439
rect 258 287 337 312
rect 266 166 322 263
rect 266 40 322 137
rect 346 40 402 137
<< ntransistor >>
rect 112 4240 152 4242
rect 184 4240 224 4242
rect 442 4240 482 4242
rect 514 4240 554 4242
rect 112 4201 152 4203
rect 184 4201 224 4203
rect 442 4201 482 4203
rect 514 4201 554 4203
rect 228 4129 248 4131
rect 185 4064 225 4066
rect 185 4025 225 4027
rect 185 3938 225 3940
rect 443 3938 483 3940
rect 185 3899 225 3901
rect 443 3899 483 3901
rect 1140 3621 1160 3623
rect 1097 3546 1137 3548
rect 1951 3546 1953 3586
rect 1990 3546 1992 3586
rect 1097 3507 1137 3509
rect 112 3283 152 3285
rect 184 3283 224 3285
rect 442 3283 482 3285
rect 514 3283 554 3285
rect 1140 3448 1160 3450
rect 1097 3381 1137 3383
rect 1097 3342 1137 3344
rect 1141 3288 1161 3290
rect 112 3244 152 3246
rect 184 3244 224 3246
rect 442 3244 482 3246
rect 514 3244 554 3246
rect 228 3172 248 3174
rect 185 3107 225 3109
rect 185 3068 225 3070
rect 757 3188 759 3228
rect 796 3188 798 3228
rect 881 3189 883 3229
rect 920 3189 922 3229
rect 996 3189 998 3229
rect 1035 3189 1037 3229
rect 1827 3289 1829 3329
rect 1866 3289 1868 3329
rect 1951 3288 1953 3328
rect 1990 3288 1992 3328
rect 2250 3783 2252 3823
rect 2289 3783 2291 3823
rect 2250 3711 2252 3751
rect 2289 3711 2291 3751
rect 2552 3712 2554 3752
rect 2591 3712 2593 3752
rect 2361 3497 2363 3517
rect 2250 3453 2252 3493
rect 2289 3453 2291 3493
rect 2426 3454 2428 3494
rect 2465 3454 2467 3494
rect 2250 3381 2252 3421
rect 2289 3381 2291 3421
rect 2552 3454 2554 3494
rect 2591 3454 2593 3494
rect 2066 3288 2068 3328
rect 2105 3288 2107 3328
rect 1106 3160 1146 3162
rect 1106 3121 1146 3123
rect 185 2981 225 2983
rect 443 2981 483 2983
rect 185 2942 225 2944
rect 443 2942 483 2944
rect 112 2804 152 2806
rect 184 2804 224 2806
rect 442 2804 482 2806
rect 514 2804 554 2806
rect 112 2765 152 2767
rect 184 2765 224 2767
rect 442 2765 482 2767
rect 514 2765 554 2767
rect 228 2693 248 2695
rect 185 2628 225 2630
rect 185 2589 225 2591
rect 881 2931 883 2971
rect 920 2931 922 2971
rect 811 2865 851 2867
rect 811 2826 851 2828
rect 787 2772 807 2774
rect 1150 3067 1170 3069
rect 1827 3068 1829 3108
rect 1866 3068 1868 3108
rect 1951 3069 1953 3109
rect 1990 3069 1992 3109
rect 2066 3069 2068 3109
rect 2105 3069 2107 3109
rect 1107 2955 1147 2957
rect 1107 2916 1147 2918
rect 1151 2862 1171 2864
rect 1151 2781 1171 2783
rect 185 2502 225 2504
rect 443 2502 483 2504
rect 185 2463 225 2465
rect 443 2463 483 2465
rect 112 2325 152 2327
rect 184 2325 224 2327
rect 442 2325 482 2327
rect 514 2325 554 2327
rect 112 2286 152 2288
rect 184 2286 224 2288
rect 442 2286 482 2288
rect 514 2286 554 2288
rect 228 2214 248 2216
rect 185 2149 225 2151
rect 185 2110 225 2112
rect 1108 2706 1148 2708
rect 1108 2667 1148 2669
rect 787 2643 807 2645
rect 1151 2608 1171 2610
rect 811 2589 851 2591
rect 811 2550 851 2552
rect 881 2446 883 2486
rect 920 2446 922 2486
rect 757 2189 759 2229
rect 796 2189 798 2229
rect 185 2023 225 2025
rect 443 2023 483 2025
rect 185 1984 225 1986
rect 443 1984 483 1986
rect 112 1846 152 1848
rect 184 1846 224 1848
rect 442 1846 482 1848
rect 514 1846 554 1848
rect 112 1807 152 1809
rect 184 1807 224 1809
rect 442 1807 482 1809
rect 514 1807 554 1809
rect 1204 2232 1206 2252
rect 881 2188 883 2228
rect 920 2188 922 2228
rect 996 2188 998 2228
rect 1035 2188 1037 2228
rect 1111 2188 1113 2228
rect 1150 2188 1152 2228
rect 1951 2811 1953 2851
rect 1990 2811 1992 2851
rect 1387 2731 1407 2733
rect 2250 3123 2252 3163
rect 2289 3123 2291 3163
rect 2250 3051 2252 3091
rect 2289 3051 2291 3091
rect 2552 3052 2554 3092
rect 2591 3052 2593 3092
rect 2361 2837 2363 2857
rect 2250 2793 2252 2833
rect 2289 2793 2291 2833
rect 2426 2794 2428 2834
rect 2465 2794 2467 2834
rect 2250 2721 2252 2761
rect 2289 2721 2291 2761
rect 2552 2794 2554 2834
rect 2591 2794 2593 2834
rect 1410 2656 1450 2658
rect 1410 2617 1450 2619
rect 1387 2558 1407 2560
rect 228 1735 248 1737
rect 185 1670 225 1672
rect 185 1631 225 1633
rect 1111 2116 1113 2156
rect 1150 2116 1152 2156
rect 757 2062 759 2102
rect 796 2062 798 2102
rect 881 2063 883 2103
rect 920 2063 922 2103
rect 996 2063 998 2103
rect 1035 2063 1037 2103
rect 1204 2092 1206 2112
rect 185 1544 225 1546
rect 443 1544 483 1546
rect 185 1505 225 1507
rect 443 1505 483 1507
rect 112 1367 152 1369
rect 184 1367 224 1369
rect 442 1367 482 1369
rect 514 1367 554 1369
rect 112 1328 152 1330
rect 184 1328 224 1330
rect 442 1328 482 1330
rect 514 1328 554 1330
rect 228 1256 248 1258
rect 185 1191 225 1193
rect 185 1152 225 1154
rect 881 1805 883 1845
rect 920 1805 922 1845
rect 811 1739 851 1741
rect 811 1700 851 1702
rect 787 1646 807 1648
rect 185 1065 225 1067
rect 443 1065 483 1067
rect 185 1026 225 1028
rect 443 1026 483 1028
rect 112 888 152 890
rect 184 888 224 890
rect 442 888 482 890
rect 514 888 554 890
rect 112 849 152 851
rect 184 849 224 851
rect 442 849 482 851
rect 514 849 554 851
rect 228 777 248 779
rect 185 712 225 714
rect 185 673 225 675
rect 185 586 225 588
rect 443 586 483 588
rect 185 547 225 549
rect 443 547 483 549
rect 112 409 152 411
rect 184 409 224 411
rect 442 409 482 411
rect 514 409 554 411
rect 112 370 152 372
rect 184 370 224 372
rect 442 370 482 372
rect 514 370 554 372
rect 228 298 248 300
rect 185 233 225 235
rect 185 194 225 196
rect 1951 2420 1953 2460
rect 1990 2420 1992 2460
rect 1450 2376 1470 2378
rect 1473 2301 1513 2303
rect 1473 2262 1513 2264
rect 1602 2206 1622 2208
rect 1450 2203 1470 2205
rect 1454 2141 1474 2143
rect 1559 2131 1599 2133
rect 1559 2092 1599 2094
rect 1477 2066 1517 2068
rect 1827 2163 1829 2203
rect 1866 2163 1868 2203
rect 1951 2162 1953 2202
rect 1990 2162 1992 2202
rect 2066 2162 2068 2202
rect 2105 2162 2107 2202
rect 1602 2033 1622 2035
rect 1477 2027 1517 2029
rect 1204 1886 1206 1906
rect 1111 1842 1113 1882
rect 1150 1842 1152 1882
rect 2250 2463 2252 2503
rect 2289 2463 2291 2503
rect 2250 2391 2252 2431
rect 2289 2391 2291 2431
rect 2552 2392 2554 2432
rect 2591 2392 2593 2432
rect 2361 2177 2363 2197
rect 2250 2133 2252 2173
rect 2289 2133 2291 2173
rect 2426 2134 2428 2174
rect 2465 2134 2467 2174
rect 2250 2061 2252 2101
rect 2289 2061 2291 2101
rect 2552 2134 2554 2174
rect 2591 2134 2593 2174
rect 1454 1968 1474 1970
rect 1108 1733 1110 1773
rect 1147 1733 1149 1773
rect 1201 1709 1203 1729
rect 1827 1942 1829 1982
rect 1866 1942 1868 1982
rect 1951 1943 1953 1983
rect 1990 1943 1992 1983
rect 2066 1943 2068 1983
rect 2105 1943 2107 1983
rect 1104 1532 1106 1572
rect 1143 1532 1145 1572
rect 1197 1508 1199 1528
rect 1197 1304 1199 1324
rect 1104 1260 1106 1300
rect 1143 1260 1145 1300
rect 1104 1159 1106 1199
rect 1143 1159 1145 1199
rect 1197 1135 1199 1155
rect 1951 1685 1953 1725
rect 1990 1685 1992 1725
rect 1547 1605 1567 1607
rect 1570 1530 1610 1532
rect 1570 1491 1610 1493
rect 1699 1435 1719 1437
rect 1547 1432 1567 1434
rect 1551 1370 1571 1372
rect 1656 1360 1696 1362
rect 1656 1321 1696 1323
rect 1574 1295 1614 1297
rect 1699 1262 1719 1264
rect 1574 1256 1614 1258
rect 2250 1803 2252 1843
rect 2289 1803 2291 1843
rect 2250 1731 2252 1771
rect 2289 1731 2291 1771
rect 2552 1732 2554 1772
rect 2591 1732 2593 1772
rect 2361 1517 2363 1537
rect 2250 1473 2252 1513
rect 2289 1473 2291 1513
rect 2426 1474 2428 1514
rect 2465 1474 2467 1514
rect 2250 1401 2252 1441
rect 2289 1401 2291 1441
rect 2552 1474 2554 1514
rect 2591 1474 2593 1514
rect 1551 1197 1571 1199
rect 1690 1173 1710 1175
rect 1647 1098 1687 1100
rect 1647 1059 1687 1061
rect 1690 1000 1710 1002
rect 2250 1143 2252 1183
rect 2289 1143 2291 1183
rect 2250 1071 2252 1111
rect 2289 1071 2291 1111
rect 2552 1072 2554 1112
rect 2591 1072 2593 1112
rect 2361 857 2363 877
rect 2250 813 2252 853
rect 2289 813 2291 853
rect 2426 814 2428 854
rect 2465 814 2467 854
rect 2250 741 2252 781
rect 2289 741 2291 781
rect 2552 814 2554 854
rect 2591 814 2593 854
rect 185 107 225 109
rect 443 107 483 109
rect 185 68 225 70
rect 443 68 483 70
<< ptransistor >>
rect 24 4240 64 4242
rect 272 4240 312 4242
rect 354 4240 394 4242
rect 602 4240 642 4242
rect 24 4201 64 4203
rect 272 4201 312 4203
rect 354 4201 394 4203
rect 602 4201 642 4203
rect 270 4129 320 4131
rect 273 4064 313 4066
rect 273 4025 313 4027
rect 273 3938 313 3940
rect 355 3938 395 3940
rect 273 3899 313 3901
rect 355 3899 395 3901
rect 2250 3871 2252 3911
rect 2289 3871 2291 3911
rect 1182 3621 1232 3623
rect 1185 3546 1225 3548
rect 1185 3507 1225 3509
rect 24 3283 64 3285
rect 272 3283 312 3285
rect 354 3283 394 3285
rect 602 3283 642 3285
rect 1182 3448 1232 3450
rect 1951 3458 1953 3498
rect 1990 3458 1992 3498
rect 1185 3381 1225 3383
rect 1827 3377 1829 3417
rect 1866 3377 1868 3417
rect 1185 3342 1225 3344
rect 1183 3288 1233 3290
rect 24 3244 64 3246
rect 272 3244 312 3246
rect 354 3244 394 3246
rect 602 3244 642 3246
rect 270 3172 320 3174
rect 273 3107 313 3109
rect 273 3068 313 3070
rect 1951 3376 1953 3416
rect 1990 3376 1992 3416
rect 2066 3376 2068 3416
rect 2105 3376 2107 3416
rect 2250 3623 2252 3663
rect 2289 3623 2291 3663
rect 2552 3624 2554 3664
rect 2591 3624 2593 3664
rect 2250 3541 2252 3581
rect 2289 3541 2291 3581
rect 2361 3539 2363 3589
rect 2426 3542 2428 3582
rect 2465 3542 2467 3582
rect 2552 3542 2554 3582
rect 2591 3542 2593 3582
rect 2250 3293 2252 3333
rect 2289 3293 2291 3333
rect 2250 3211 2252 3251
rect 2289 3211 2291 3251
rect 757 3100 759 3140
rect 796 3100 798 3140
rect 1194 3160 1234 3162
rect 881 3101 883 3141
rect 920 3101 922 3141
rect 996 3101 998 3141
rect 1035 3101 1037 3141
rect 1194 3121 1234 3123
rect 881 3019 883 3059
rect 920 3019 922 3059
rect 273 2981 313 2983
rect 355 2981 395 2983
rect 273 2942 313 2944
rect 355 2942 395 2944
rect 24 2804 64 2806
rect 272 2804 312 2806
rect 354 2804 394 2806
rect 602 2804 642 2806
rect 24 2765 64 2767
rect 272 2765 312 2767
rect 354 2765 394 2767
rect 602 2765 642 2767
rect 270 2693 320 2695
rect 273 2628 313 2630
rect 273 2589 313 2591
rect 723 2865 763 2867
rect 723 2826 763 2828
rect 715 2772 765 2774
rect 1192 3067 1242 3069
rect 1827 2980 1829 3020
rect 1866 2980 1868 3020
rect 1195 2955 1235 2957
rect 1195 2916 1235 2918
rect 1951 2981 1953 3021
rect 1990 2981 1992 3021
rect 2066 2981 2068 3021
rect 2105 2981 2107 3021
rect 1951 2899 1953 2939
rect 1990 2899 1992 2939
rect 1193 2862 1243 2864
rect 1193 2781 1243 2783
rect 273 2502 313 2504
rect 355 2502 395 2504
rect 273 2463 313 2465
rect 355 2463 395 2465
rect 24 2325 64 2327
rect 272 2325 312 2327
rect 354 2325 394 2327
rect 602 2325 642 2327
rect 24 2286 64 2288
rect 272 2286 312 2288
rect 354 2286 394 2288
rect 602 2286 642 2288
rect 270 2214 320 2216
rect 273 2149 313 2151
rect 273 2110 313 2112
rect 1196 2706 1236 2708
rect 1196 2667 1236 2669
rect 715 2643 765 2645
rect 1193 2608 1243 2610
rect 723 2589 763 2591
rect 723 2550 763 2552
rect 757 2277 759 2317
rect 796 2277 798 2317
rect 881 2358 883 2398
rect 920 2358 922 2398
rect 881 2276 883 2316
rect 920 2276 922 2316
rect 996 2276 998 2316
rect 1035 2276 1037 2316
rect 1111 2276 1113 2316
rect 1150 2276 1152 2316
rect 273 2023 313 2025
rect 355 2023 395 2025
rect 273 1984 313 1986
rect 355 1984 395 1986
rect 24 1846 64 1848
rect 272 1846 312 1848
rect 354 1846 394 1848
rect 602 1846 642 1848
rect 24 1807 64 1809
rect 272 1807 312 1809
rect 354 1807 394 1809
rect 602 1807 642 1809
rect 1204 2274 1206 2324
rect 1315 2731 1365 2733
rect 2250 2963 2252 3003
rect 2289 2963 2291 3003
rect 2552 2964 2554 3004
rect 2591 2964 2593 3004
rect 2250 2881 2252 2921
rect 2289 2881 2291 2921
rect 2361 2879 2363 2929
rect 2426 2882 2428 2922
rect 2465 2882 2467 2922
rect 2552 2882 2554 2922
rect 2591 2882 2593 2922
rect 1322 2656 1362 2658
rect 2250 2633 2252 2673
rect 2289 2633 2291 2673
rect 1322 2617 1362 2619
rect 1315 2558 1365 2560
rect 270 1735 320 1737
rect 273 1670 313 1672
rect 273 1631 313 1633
rect 757 1974 759 2014
rect 796 1974 798 2014
rect 881 1975 883 2015
rect 920 1975 922 2015
rect 996 1975 998 2015
rect 1035 1975 1037 2015
rect 881 1893 883 1933
rect 920 1893 922 1933
rect 273 1544 313 1546
rect 355 1544 395 1546
rect 273 1505 313 1507
rect 355 1505 395 1507
rect 24 1367 64 1369
rect 272 1367 312 1369
rect 354 1367 394 1369
rect 602 1367 642 1369
rect 24 1328 64 1330
rect 272 1328 312 1330
rect 354 1328 394 1330
rect 602 1328 642 1330
rect 270 1256 320 1258
rect 273 1191 313 1193
rect 273 1152 313 1154
rect 723 1739 763 1741
rect 723 1700 763 1702
rect 715 1646 765 1648
rect 273 1065 313 1067
rect 355 1065 395 1067
rect 273 1026 313 1028
rect 355 1026 395 1028
rect 24 888 64 890
rect 272 888 312 890
rect 354 888 394 890
rect 602 888 642 890
rect 24 849 64 851
rect 272 849 312 851
rect 354 849 394 851
rect 602 849 642 851
rect 270 777 320 779
rect 273 712 313 714
rect 273 673 313 675
rect 273 586 313 588
rect 355 586 395 588
rect 273 547 313 549
rect 355 547 395 549
rect 24 409 64 411
rect 272 409 312 411
rect 354 409 394 411
rect 602 409 642 411
rect 24 370 64 372
rect 272 370 312 372
rect 354 370 394 372
rect 602 370 642 372
rect 270 298 320 300
rect 273 233 313 235
rect 273 194 313 196
rect 1111 2028 1113 2068
rect 1150 2028 1152 2068
rect 1204 2020 1206 2070
rect 2250 2551 2252 2591
rect 2289 2551 2291 2591
rect 1378 2376 1428 2378
rect 1951 2332 1953 2372
rect 1990 2332 1992 2372
rect 1385 2301 1425 2303
rect 1385 2262 1425 2264
rect 1827 2251 1829 2291
rect 1866 2251 1868 2291
rect 1644 2206 1694 2208
rect 1378 2203 1428 2205
rect 1951 2250 1953 2290
rect 1990 2250 1992 2290
rect 1382 2141 1432 2143
rect 1647 2131 1687 2133
rect 1647 2092 1687 2094
rect 1389 2066 1429 2068
rect 2066 2250 2068 2290
rect 2105 2250 2107 2290
rect 1644 2033 1694 2035
rect 1389 2027 1429 2029
rect 1111 1930 1113 1970
rect 1150 1930 1152 1970
rect 1204 1928 1206 1978
rect 2250 2303 2252 2343
rect 2289 2303 2291 2343
rect 2552 2304 2554 2344
rect 2591 2304 2593 2344
rect 2250 2221 2252 2261
rect 2289 2221 2291 2261
rect 2361 2219 2363 2269
rect 2426 2222 2428 2262
rect 2465 2222 2467 2262
rect 2552 2222 2554 2262
rect 2591 2222 2593 2262
rect 1382 1968 1432 1970
rect 1108 1645 1110 1685
rect 1147 1645 1149 1685
rect 1201 1637 1203 1687
rect 2250 1973 2252 2013
rect 2289 1973 2291 2013
rect 1104 1444 1106 1484
rect 1143 1444 1145 1484
rect 1197 1436 1199 1486
rect 1104 1348 1106 1388
rect 1143 1348 1145 1388
rect 1197 1346 1199 1396
rect 1104 1071 1106 1111
rect 1143 1071 1145 1111
rect 1197 1063 1199 1113
rect 1827 1854 1829 1894
rect 1866 1854 1868 1894
rect 1951 1855 1953 1895
rect 1990 1855 1992 1895
rect 2066 1855 2068 1895
rect 2105 1855 2107 1895
rect 1951 1773 1953 1813
rect 1990 1773 1992 1813
rect 1475 1605 1525 1607
rect 1482 1530 1522 1532
rect 1482 1491 1522 1493
rect 1741 1435 1791 1437
rect 1475 1432 1525 1434
rect 1479 1370 1529 1372
rect 1744 1360 1784 1362
rect 1744 1321 1784 1323
rect 1486 1295 1526 1297
rect 1741 1262 1791 1264
rect 1486 1256 1526 1258
rect 2250 1891 2252 1931
rect 2289 1891 2291 1931
rect 2250 1643 2252 1683
rect 2289 1643 2291 1683
rect 2552 1644 2554 1684
rect 2591 1644 2593 1684
rect 2250 1561 2252 1601
rect 2289 1561 2291 1601
rect 2361 1559 2363 1609
rect 2426 1562 2428 1602
rect 2465 1562 2467 1602
rect 2552 1562 2554 1602
rect 2591 1562 2593 1602
rect 2250 1313 2252 1353
rect 2289 1313 2291 1353
rect 2250 1231 2252 1271
rect 2289 1231 2291 1271
rect 1479 1197 1529 1199
rect 1732 1173 1782 1175
rect 1735 1098 1775 1100
rect 1735 1059 1775 1061
rect 1732 1000 1782 1002
rect 2250 983 2252 1023
rect 2289 983 2291 1023
rect 2552 984 2554 1024
rect 2591 984 2593 1024
rect 2250 901 2252 941
rect 2289 901 2291 941
rect 2361 899 2363 949
rect 2426 902 2428 942
rect 2465 902 2467 942
rect 2552 902 2554 942
rect 2591 902 2593 942
rect 2250 653 2252 693
rect 2289 653 2291 693
rect 273 107 313 109
rect 355 107 395 109
rect 273 68 313 70
rect 355 68 395 70
<< ndiffusion >>
rect 112 4259 152 4262
rect 150 4252 152 4259
rect 112 4242 152 4252
rect 184 4259 224 4262
rect 184 4252 186 4259
rect 184 4242 224 4252
rect 112 4203 152 4240
rect 184 4203 224 4240
rect 442 4259 482 4262
rect 480 4252 482 4259
rect 442 4242 482 4252
rect 514 4259 554 4262
rect 514 4252 516 4259
rect 514 4242 554 4252
rect 442 4203 482 4240
rect 514 4203 554 4240
rect 112 4193 152 4201
rect 150 4186 152 4193
rect 112 4182 152 4186
rect 184 4193 224 4201
rect 184 4186 186 4193
rect 184 4182 224 4186
rect 442 4193 482 4201
rect 480 4186 482 4193
rect 442 4182 482 4186
rect 514 4193 554 4201
rect 514 4186 516 4193
rect 514 4182 554 4186
rect 228 4131 248 4132
rect 228 4128 248 4129
rect 185 4083 225 4086
rect 185 4076 187 4083
rect 185 4066 225 4076
rect 185 4027 225 4064
rect 185 4017 225 4025
rect 185 4010 187 4017
rect 185 4006 225 4010
rect 185 3957 225 3960
rect 185 3950 187 3957
rect 185 3940 225 3950
rect 443 3957 483 3960
rect 185 3901 225 3938
rect 481 3950 483 3957
rect 443 3940 483 3950
rect 443 3901 483 3938
rect 185 3891 225 3899
rect 185 3884 187 3891
rect 185 3880 225 3884
rect 443 3891 483 3899
rect 481 3884 483 3891
rect 443 3880 483 3884
rect 1140 3623 1160 3624
rect 1140 3620 1160 3621
rect 1097 3565 1137 3568
rect 1097 3558 1099 3565
rect 1097 3548 1137 3558
rect 1097 3509 1137 3546
rect 1931 3584 1951 3586
rect 1931 3546 1934 3584
rect 1941 3546 1951 3584
rect 1953 3546 1990 3586
rect 1992 3584 2011 3586
rect 1992 3546 2000 3584
rect 2007 3546 2011 3584
rect 1097 3499 1137 3507
rect 112 3302 152 3305
rect 150 3295 152 3302
rect 112 3285 152 3295
rect 184 3302 224 3305
rect 184 3295 186 3302
rect 184 3285 224 3295
rect 112 3246 152 3283
rect 184 3246 224 3283
rect 442 3302 482 3305
rect 480 3295 482 3302
rect 442 3285 482 3295
rect 514 3302 554 3305
rect 514 3295 516 3302
rect 514 3285 554 3295
rect 442 3246 482 3283
rect 514 3246 554 3283
rect 1097 3492 1099 3499
rect 1097 3488 1137 3492
rect 1140 3450 1160 3451
rect 1140 3447 1160 3448
rect 1097 3400 1137 3403
rect 1097 3393 1099 3400
rect 1097 3383 1137 3393
rect 1097 3344 1137 3381
rect 1097 3334 1137 3342
rect 1097 3327 1099 3334
rect 1097 3323 1137 3327
rect 1141 3290 1161 3291
rect 1141 3287 1161 3288
rect 112 3236 152 3244
rect 150 3229 152 3236
rect 112 3225 152 3229
rect 184 3236 224 3244
rect 184 3229 186 3236
rect 184 3225 224 3229
rect 442 3236 482 3244
rect 480 3229 482 3236
rect 442 3225 482 3229
rect 514 3236 554 3244
rect 514 3229 516 3236
rect 514 3225 554 3229
rect 228 3174 248 3175
rect 228 3171 248 3172
rect 185 3126 225 3129
rect 185 3119 187 3126
rect 185 3109 225 3119
rect 185 3070 225 3107
rect 185 3060 225 3068
rect 185 3053 187 3060
rect 185 3049 225 3053
rect 737 3226 757 3228
rect 737 3188 740 3226
rect 747 3188 757 3226
rect 759 3188 796 3228
rect 798 3226 817 3228
rect 798 3188 806 3226
rect 813 3188 817 3226
rect 861 3227 881 3229
rect 861 3189 864 3227
rect 871 3189 881 3227
rect 883 3189 920 3229
rect 922 3227 941 3229
rect 922 3189 930 3227
rect 937 3189 941 3227
rect 976 3227 996 3229
rect 976 3189 979 3227
rect 986 3189 996 3227
rect 998 3189 1035 3229
rect 1037 3227 1056 3229
rect 1037 3189 1045 3227
rect 1052 3189 1056 3227
rect 1807 3291 1810 3329
rect 1817 3291 1827 3329
rect 1807 3289 1827 3291
rect 1829 3289 1866 3329
rect 1868 3291 1876 3329
rect 1883 3291 1887 3329
rect 1868 3289 1887 3291
rect 1931 3290 1934 3328
rect 1941 3290 1951 3328
rect 1931 3288 1951 3290
rect 1953 3288 1990 3328
rect 1992 3290 2000 3328
rect 2007 3290 2011 3328
rect 1992 3288 2011 3290
rect 2230 3785 2233 3823
rect 2240 3785 2250 3823
rect 2230 3783 2250 3785
rect 2252 3783 2289 3823
rect 2291 3785 2299 3823
rect 2306 3785 2310 3823
rect 2291 3783 2310 3785
rect 2230 3749 2250 3751
rect 2230 3711 2233 3749
rect 2240 3711 2250 3749
rect 2252 3711 2289 3751
rect 2291 3749 2310 3751
rect 2291 3711 2299 3749
rect 2306 3711 2310 3749
rect 2532 3750 2552 3752
rect 2532 3712 2535 3750
rect 2542 3712 2552 3750
rect 2554 3712 2591 3752
rect 2593 3750 2612 3752
rect 2593 3712 2601 3750
rect 2608 3712 2612 3750
rect 2360 3497 2361 3517
rect 2363 3497 2364 3517
rect 2230 3455 2233 3493
rect 2240 3455 2250 3493
rect 2230 3453 2250 3455
rect 2252 3453 2289 3493
rect 2291 3455 2299 3493
rect 2306 3455 2310 3493
rect 2291 3453 2310 3455
rect 2406 3456 2409 3494
rect 2416 3456 2426 3494
rect 2406 3454 2426 3456
rect 2428 3454 2465 3494
rect 2467 3456 2475 3494
rect 2482 3456 2486 3494
rect 2467 3454 2486 3456
rect 2230 3419 2250 3421
rect 2230 3381 2233 3419
rect 2240 3381 2250 3419
rect 2252 3381 2289 3421
rect 2291 3419 2310 3421
rect 2291 3381 2299 3419
rect 2306 3381 2310 3419
rect 2532 3456 2535 3494
rect 2542 3456 2552 3494
rect 2532 3454 2552 3456
rect 2554 3454 2591 3494
rect 2593 3456 2601 3494
rect 2608 3456 2612 3494
rect 2593 3454 2612 3456
rect 2046 3290 2049 3328
rect 2056 3290 2066 3328
rect 2046 3288 2066 3290
rect 2068 3288 2105 3328
rect 2107 3290 2115 3328
rect 2122 3290 2126 3328
rect 2107 3288 2126 3290
rect 1106 3179 1146 3182
rect 1106 3172 1108 3179
rect 1106 3162 1146 3172
rect 1106 3123 1146 3160
rect 185 3000 225 3003
rect 185 2993 187 3000
rect 185 2983 225 2993
rect 443 3000 483 3003
rect 185 2944 225 2981
rect 481 2993 483 3000
rect 443 2983 483 2993
rect 443 2944 483 2981
rect 185 2934 225 2942
rect 185 2927 187 2934
rect 185 2923 225 2927
rect 443 2934 483 2942
rect 481 2927 483 2934
rect 443 2923 483 2927
rect 112 2823 152 2826
rect 150 2816 152 2823
rect 112 2806 152 2816
rect 184 2823 224 2826
rect 184 2816 186 2823
rect 184 2806 224 2816
rect 112 2767 152 2804
rect 184 2767 224 2804
rect 442 2823 482 2826
rect 480 2816 482 2823
rect 442 2806 482 2816
rect 514 2823 554 2826
rect 514 2816 516 2823
rect 514 2806 554 2816
rect 442 2767 482 2804
rect 514 2767 554 2804
rect 112 2757 152 2765
rect 150 2750 152 2757
rect 112 2746 152 2750
rect 184 2757 224 2765
rect 184 2750 186 2757
rect 184 2746 224 2750
rect 442 2757 482 2765
rect 480 2750 482 2757
rect 442 2746 482 2750
rect 514 2757 554 2765
rect 514 2750 516 2757
rect 514 2746 554 2750
rect 228 2695 248 2696
rect 228 2692 248 2693
rect 185 2647 225 2650
rect 185 2640 187 2647
rect 185 2630 225 2640
rect 185 2591 225 2628
rect 185 2581 225 2589
rect 185 2574 187 2581
rect 185 2570 225 2574
rect 861 2933 864 2971
rect 871 2933 881 2971
rect 861 2931 881 2933
rect 883 2931 920 2971
rect 922 2933 930 2971
rect 937 2933 941 2971
rect 922 2931 941 2933
rect 811 2884 851 2887
rect 849 2877 851 2884
rect 811 2867 851 2877
rect 811 2828 851 2865
rect 811 2818 851 2826
rect 849 2811 851 2818
rect 811 2807 851 2811
rect 787 2774 807 2775
rect 787 2771 807 2772
rect 1106 3113 1146 3121
rect 1106 3106 1108 3113
rect 1106 3102 1146 3106
rect 1807 3106 1827 3108
rect 1150 3069 1170 3070
rect 1807 3068 1810 3106
rect 1817 3068 1827 3106
rect 1829 3068 1866 3108
rect 1868 3106 1887 3108
rect 1868 3068 1876 3106
rect 1883 3068 1887 3106
rect 1931 3107 1951 3109
rect 1931 3069 1934 3107
rect 1941 3069 1951 3107
rect 1953 3069 1990 3109
rect 1992 3107 2011 3109
rect 1992 3069 2000 3107
rect 2007 3069 2011 3107
rect 2046 3107 2066 3109
rect 2046 3069 2049 3107
rect 2056 3069 2066 3107
rect 2068 3069 2105 3109
rect 2107 3107 2126 3109
rect 2107 3069 2115 3107
rect 2122 3069 2126 3107
rect 1150 3066 1170 3067
rect 1107 2974 1147 2977
rect 1107 2967 1109 2974
rect 1107 2957 1147 2967
rect 1107 2918 1147 2955
rect 1107 2908 1147 2916
rect 1107 2901 1109 2908
rect 1107 2897 1147 2901
rect 1151 2864 1171 2865
rect 1151 2861 1171 2862
rect 1151 2783 1171 2784
rect 1151 2780 1171 2781
rect 185 2521 225 2524
rect 185 2514 187 2521
rect 185 2504 225 2514
rect 443 2521 483 2524
rect 185 2465 225 2502
rect 481 2514 483 2521
rect 443 2504 483 2514
rect 443 2465 483 2502
rect 185 2455 225 2463
rect 185 2448 187 2455
rect 185 2444 225 2448
rect 443 2455 483 2463
rect 481 2448 483 2455
rect 443 2444 483 2448
rect 112 2344 152 2347
rect 150 2337 152 2344
rect 112 2327 152 2337
rect 184 2344 224 2347
rect 184 2337 186 2344
rect 184 2327 224 2337
rect 112 2288 152 2325
rect 184 2288 224 2325
rect 442 2344 482 2347
rect 480 2337 482 2344
rect 442 2327 482 2337
rect 514 2344 554 2347
rect 514 2337 516 2344
rect 514 2327 554 2337
rect 442 2288 482 2325
rect 514 2288 554 2325
rect 112 2278 152 2286
rect 150 2271 152 2278
rect 112 2267 152 2271
rect 184 2278 224 2286
rect 184 2271 186 2278
rect 184 2267 224 2271
rect 442 2278 482 2286
rect 480 2271 482 2278
rect 442 2267 482 2271
rect 514 2278 554 2286
rect 514 2271 516 2278
rect 514 2267 554 2271
rect 228 2216 248 2217
rect 228 2213 248 2214
rect 185 2168 225 2171
rect 185 2161 187 2168
rect 185 2151 225 2161
rect 185 2112 225 2149
rect 185 2102 225 2110
rect 185 2095 187 2102
rect 185 2091 225 2095
rect 1108 2725 1148 2728
rect 1108 2718 1110 2725
rect 1108 2708 1148 2718
rect 1108 2669 1148 2706
rect 1108 2659 1148 2667
rect 1108 2652 1110 2659
rect 1108 2648 1148 2652
rect 787 2645 807 2646
rect 787 2642 807 2643
rect 1151 2610 1171 2611
rect 811 2606 851 2610
rect 849 2599 851 2606
rect 1151 2607 1171 2608
rect 811 2591 851 2599
rect 811 2552 851 2589
rect 811 2540 851 2550
rect 849 2533 851 2540
rect 811 2530 851 2533
rect 861 2484 881 2486
rect 861 2446 864 2484
rect 871 2446 881 2484
rect 883 2446 920 2486
rect 922 2484 941 2486
rect 922 2446 930 2484
rect 937 2446 941 2484
rect 737 2191 740 2229
rect 747 2191 757 2229
rect 737 2189 757 2191
rect 759 2189 796 2229
rect 798 2191 806 2229
rect 813 2191 817 2229
rect 798 2189 817 2191
rect 185 2042 225 2045
rect 185 2035 187 2042
rect 185 2025 225 2035
rect 443 2042 483 2045
rect 185 1986 225 2023
rect 481 2035 483 2042
rect 443 2025 483 2035
rect 443 1986 483 2023
rect 185 1976 225 1984
rect 185 1969 187 1976
rect 185 1965 225 1969
rect 443 1976 483 1984
rect 481 1969 483 1976
rect 443 1965 483 1969
rect 112 1865 152 1868
rect 150 1858 152 1865
rect 112 1848 152 1858
rect 184 1865 224 1868
rect 184 1858 186 1865
rect 184 1848 224 1858
rect 112 1809 152 1846
rect 184 1809 224 1846
rect 442 1865 482 1868
rect 480 1858 482 1865
rect 442 1848 482 1858
rect 514 1865 554 1868
rect 514 1858 516 1865
rect 514 1848 554 1858
rect 442 1809 482 1846
rect 514 1809 554 1846
rect 112 1799 152 1807
rect 150 1792 152 1799
rect 112 1788 152 1792
rect 184 1799 224 1807
rect 184 1792 186 1799
rect 184 1788 224 1792
rect 442 1799 482 1807
rect 480 1792 482 1799
rect 442 1788 482 1792
rect 514 1799 554 1807
rect 514 1792 516 1799
rect 514 1788 554 1792
rect 1203 2232 1204 2252
rect 1206 2232 1207 2252
rect 861 2190 864 2228
rect 871 2190 881 2228
rect 861 2188 881 2190
rect 883 2188 920 2228
rect 922 2190 930 2228
rect 937 2190 941 2228
rect 922 2188 941 2190
rect 976 2190 979 2228
rect 986 2190 996 2228
rect 976 2188 996 2190
rect 998 2188 1035 2228
rect 1037 2190 1045 2228
rect 1052 2190 1056 2228
rect 1037 2188 1056 2190
rect 1091 2190 1094 2228
rect 1101 2190 1111 2228
rect 1091 2188 1111 2190
rect 1113 2188 1150 2228
rect 1152 2190 1160 2228
rect 1167 2190 1171 2228
rect 1152 2188 1171 2190
rect 1931 2813 1934 2851
rect 1941 2813 1951 2851
rect 1931 2811 1951 2813
rect 1953 2811 1990 2851
rect 1992 2813 2000 2851
rect 2007 2813 2011 2851
rect 1992 2811 2011 2813
rect 1387 2733 1407 2734
rect 1387 2730 1407 2731
rect 2230 3125 2233 3163
rect 2240 3125 2250 3163
rect 2230 3123 2250 3125
rect 2252 3123 2289 3163
rect 2291 3125 2299 3163
rect 2306 3125 2310 3163
rect 2291 3123 2310 3125
rect 2230 3089 2250 3091
rect 2230 3051 2233 3089
rect 2240 3051 2250 3089
rect 2252 3051 2289 3091
rect 2291 3089 2310 3091
rect 2291 3051 2299 3089
rect 2306 3051 2310 3089
rect 2532 3090 2552 3092
rect 2532 3052 2535 3090
rect 2542 3052 2552 3090
rect 2554 3052 2591 3092
rect 2593 3090 2612 3092
rect 2593 3052 2601 3090
rect 2608 3052 2612 3090
rect 2360 2837 2361 2857
rect 2363 2837 2364 2857
rect 2230 2795 2233 2833
rect 2240 2795 2250 2833
rect 2230 2793 2250 2795
rect 2252 2793 2289 2833
rect 2291 2795 2299 2833
rect 2306 2795 2310 2833
rect 2291 2793 2310 2795
rect 2406 2796 2409 2834
rect 2416 2796 2426 2834
rect 2406 2794 2426 2796
rect 2428 2794 2465 2834
rect 2467 2796 2475 2834
rect 2482 2796 2486 2834
rect 2467 2794 2486 2796
rect 2230 2759 2250 2761
rect 2230 2721 2233 2759
rect 2240 2721 2250 2759
rect 2252 2721 2289 2761
rect 2291 2759 2310 2761
rect 2291 2721 2299 2759
rect 2306 2721 2310 2759
rect 1410 2675 1450 2678
rect 1448 2668 1450 2675
rect 2532 2796 2535 2834
rect 2542 2796 2552 2834
rect 2532 2794 2552 2796
rect 2554 2794 2591 2834
rect 2593 2796 2601 2834
rect 2608 2796 2612 2834
rect 2593 2794 2612 2796
rect 1410 2658 1450 2668
rect 1410 2619 1450 2656
rect 1410 2609 1450 2617
rect 1448 2602 1450 2609
rect 1410 2598 1450 2602
rect 1387 2560 1407 2561
rect 1387 2557 1407 2558
rect 1091 2154 1111 2156
rect 228 1737 248 1738
rect 228 1734 248 1735
rect 185 1689 225 1692
rect 185 1682 187 1689
rect 185 1672 225 1682
rect 185 1633 225 1670
rect 185 1623 225 1631
rect 185 1616 187 1623
rect 185 1612 225 1616
rect 1091 2116 1094 2154
rect 1101 2116 1111 2154
rect 1113 2116 1150 2156
rect 1152 2154 1171 2156
rect 1152 2116 1160 2154
rect 1167 2116 1171 2154
rect 737 2100 757 2102
rect 737 2062 740 2100
rect 747 2062 757 2100
rect 759 2062 796 2102
rect 798 2100 817 2102
rect 798 2062 806 2100
rect 813 2062 817 2100
rect 861 2101 881 2103
rect 861 2063 864 2101
rect 871 2063 881 2101
rect 883 2063 920 2103
rect 922 2101 941 2103
rect 922 2063 930 2101
rect 937 2063 941 2101
rect 976 2101 996 2103
rect 976 2063 979 2101
rect 986 2063 996 2101
rect 998 2063 1035 2103
rect 1037 2101 1056 2103
rect 1037 2063 1045 2101
rect 1052 2063 1056 2101
rect 1203 2092 1204 2112
rect 1206 2092 1207 2112
rect 185 1563 225 1566
rect 185 1556 187 1563
rect 185 1546 225 1556
rect 443 1563 483 1566
rect 185 1507 225 1544
rect 481 1556 483 1563
rect 443 1546 483 1556
rect 443 1507 483 1544
rect 185 1497 225 1505
rect 185 1490 187 1497
rect 185 1486 225 1490
rect 443 1497 483 1505
rect 481 1490 483 1497
rect 443 1486 483 1490
rect 112 1386 152 1389
rect 150 1379 152 1386
rect 112 1369 152 1379
rect 184 1386 224 1389
rect 184 1379 186 1386
rect 184 1369 224 1379
rect 112 1330 152 1367
rect 184 1330 224 1367
rect 442 1386 482 1389
rect 480 1379 482 1386
rect 442 1369 482 1379
rect 514 1386 554 1389
rect 514 1379 516 1386
rect 514 1369 554 1379
rect 442 1330 482 1367
rect 514 1330 554 1367
rect 112 1320 152 1328
rect 150 1313 152 1320
rect 112 1309 152 1313
rect 184 1320 224 1328
rect 184 1313 186 1320
rect 184 1309 224 1313
rect 442 1320 482 1328
rect 480 1313 482 1320
rect 442 1309 482 1313
rect 514 1320 554 1328
rect 514 1313 516 1320
rect 514 1309 554 1313
rect 228 1258 248 1259
rect 228 1255 248 1256
rect 185 1210 225 1213
rect 185 1203 187 1210
rect 185 1193 225 1203
rect 185 1154 225 1191
rect 185 1144 225 1152
rect 185 1137 187 1144
rect 185 1133 225 1137
rect 861 1807 864 1845
rect 871 1807 881 1845
rect 861 1805 881 1807
rect 883 1805 920 1845
rect 922 1807 930 1845
rect 937 1807 941 1845
rect 922 1805 941 1807
rect 811 1758 851 1761
rect 849 1751 851 1758
rect 811 1741 851 1751
rect 811 1702 851 1739
rect 811 1692 851 1700
rect 849 1685 851 1692
rect 811 1681 851 1685
rect 787 1648 807 1649
rect 787 1645 807 1646
rect 185 1084 225 1087
rect 185 1077 187 1084
rect 185 1067 225 1077
rect 443 1084 483 1087
rect 185 1028 225 1065
rect 481 1077 483 1084
rect 443 1067 483 1077
rect 443 1028 483 1065
rect 185 1018 225 1026
rect 185 1011 187 1018
rect 185 1007 225 1011
rect 443 1018 483 1026
rect 481 1011 483 1018
rect 443 1007 483 1011
rect 112 907 152 910
rect 150 900 152 907
rect 112 890 152 900
rect 184 907 224 910
rect 184 900 186 907
rect 184 890 224 900
rect 112 851 152 888
rect 184 851 224 888
rect 442 907 482 910
rect 480 900 482 907
rect 442 890 482 900
rect 514 907 554 910
rect 514 900 516 907
rect 514 890 554 900
rect 442 851 482 888
rect 514 851 554 888
rect 112 841 152 849
rect 150 834 152 841
rect 112 830 152 834
rect 184 841 224 849
rect 184 834 186 841
rect 184 830 224 834
rect 442 841 482 849
rect 480 834 482 841
rect 442 830 482 834
rect 514 841 554 849
rect 514 834 516 841
rect 514 830 554 834
rect 228 779 248 780
rect 228 776 248 777
rect 185 731 225 734
rect 185 724 187 731
rect 185 714 225 724
rect 185 675 225 712
rect 185 665 225 673
rect 185 658 187 665
rect 185 654 225 658
rect 185 605 225 608
rect 185 598 187 605
rect 185 588 225 598
rect 443 605 483 608
rect 185 549 225 586
rect 481 598 483 605
rect 443 588 483 598
rect 443 549 483 586
rect 185 539 225 547
rect 185 532 187 539
rect 185 528 225 532
rect 443 539 483 547
rect 481 532 483 539
rect 443 528 483 532
rect 112 428 152 431
rect 150 421 152 428
rect 112 411 152 421
rect 184 428 224 431
rect 184 421 186 428
rect 184 411 224 421
rect 112 372 152 409
rect 184 372 224 409
rect 442 428 482 431
rect 480 421 482 428
rect 442 411 482 421
rect 514 428 554 431
rect 514 421 516 428
rect 514 411 554 421
rect 442 372 482 409
rect 514 372 554 409
rect 112 362 152 370
rect 150 355 152 362
rect 112 351 152 355
rect 184 362 224 370
rect 184 355 186 362
rect 184 351 224 355
rect 442 362 482 370
rect 480 355 482 362
rect 442 351 482 355
rect 514 362 554 370
rect 514 355 516 362
rect 514 351 554 355
rect 228 300 248 301
rect 228 297 248 298
rect 185 252 225 255
rect 185 245 187 252
rect 185 235 225 245
rect 185 196 225 233
rect 185 186 225 194
rect 185 179 187 186
rect 185 175 225 179
rect 1931 2458 1951 2460
rect 1931 2420 1934 2458
rect 1941 2420 1951 2458
rect 1953 2420 1990 2460
rect 1992 2458 2011 2460
rect 1992 2420 2000 2458
rect 2007 2420 2011 2458
rect 1450 2378 1470 2379
rect 1450 2375 1470 2376
rect 1473 2320 1513 2323
rect 1511 2313 1513 2320
rect 1473 2303 1513 2313
rect 1473 2264 1513 2301
rect 1473 2254 1513 2262
rect 1511 2247 1513 2254
rect 1473 2243 1513 2247
rect 1602 2208 1622 2209
rect 1450 2205 1470 2206
rect 1602 2205 1622 2206
rect 1450 2202 1470 2203
rect 1559 2150 1599 2153
rect 1454 2143 1474 2144
rect 1559 2143 1561 2150
rect 1454 2140 1474 2141
rect 1559 2133 1599 2143
rect 1559 2094 1599 2131
rect 1477 2085 1517 2088
rect 1515 2078 1517 2085
rect 1477 2068 1517 2078
rect 1559 2084 1599 2092
rect 1559 2077 1561 2084
rect 1559 2073 1599 2077
rect 1477 2029 1517 2066
rect 1807 2165 1810 2203
rect 1817 2165 1827 2203
rect 1807 2163 1827 2165
rect 1829 2163 1866 2203
rect 1868 2165 1876 2203
rect 1883 2165 1887 2203
rect 1868 2163 1887 2165
rect 1931 2164 1934 2202
rect 1941 2164 1951 2202
rect 1931 2162 1951 2164
rect 1953 2162 1990 2202
rect 1992 2164 2000 2202
rect 2007 2164 2011 2202
rect 1992 2162 2011 2164
rect 2046 2164 2049 2202
rect 2056 2164 2066 2202
rect 2046 2162 2066 2164
rect 2068 2162 2105 2202
rect 2107 2164 2115 2202
rect 2122 2164 2126 2202
rect 2107 2162 2126 2164
rect 1602 2035 1622 2036
rect 1602 2032 1622 2033
rect 1477 2019 1517 2027
rect 1515 2012 1517 2019
rect 1477 2008 1517 2012
rect 1203 1886 1204 1906
rect 1206 1886 1207 1906
rect 1091 1844 1094 1882
rect 1101 1844 1111 1882
rect 1091 1842 1111 1844
rect 1113 1842 1150 1882
rect 1152 1844 1160 1882
rect 1167 1844 1171 1882
rect 1152 1842 1171 1844
rect 2230 2465 2233 2503
rect 2240 2465 2250 2503
rect 2230 2463 2250 2465
rect 2252 2463 2289 2503
rect 2291 2465 2299 2503
rect 2306 2465 2310 2503
rect 2291 2463 2310 2465
rect 2230 2429 2250 2431
rect 2230 2391 2233 2429
rect 2240 2391 2250 2429
rect 2252 2391 2289 2431
rect 2291 2429 2310 2431
rect 2291 2391 2299 2429
rect 2306 2391 2310 2429
rect 2532 2430 2552 2432
rect 2532 2392 2535 2430
rect 2542 2392 2552 2430
rect 2554 2392 2591 2432
rect 2593 2430 2612 2432
rect 2593 2392 2601 2430
rect 2608 2392 2612 2430
rect 2360 2177 2361 2197
rect 2363 2177 2364 2197
rect 2230 2135 2233 2173
rect 2240 2135 2250 2173
rect 2230 2133 2250 2135
rect 2252 2133 2289 2173
rect 2291 2135 2299 2173
rect 2306 2135 2310 2173
rect 2291 2133 2310 2135
rect 2406 2136 2409 2174
rect 2416 2136 2426 2174
rect 2406 2134 2426 2136
rect 2428 2134 2465 2174
rect 2467 2136 2475 2174
rect 2482 2136 2486 2174
rect 2467 2134 2486 2136
rect 2230 2099 2250 2101
rect 2230 2061 2233 2099
rect 2240 2061 2250 2099
rect 2252 2061 2289 2101
rect 2291 2099 2310 2101
rect 2291 2061 2299 2099
rect 2306 2061 2310 2099
rect 2532 2136 2535 2174
rect 2542 2136 2552 2174
rect 2532 2134 2552 2136
rect 2554 2134 2591 2174
rect 2593 2136 2601 2174
rect 2608 2136 2612 2174
rect 2593 2134 2612 2136
rect 1807 1980 1827 1982
rect 1454 1970 1474 1971
rect 1088 1771 1108 1773
rect 1088 1733 1091 1771
rect 1098 1733 1108 1771
rect 1110 1733 1147 1773
rect 1149 1771 1168 1773
rect 1149 1733 1157 1771
rect 1164 1733 1168 1771
rect 1200 1709 1201 1729
rect 1203 1709 1204 1729
rect 1454 1967 1474 1968
rect 1807 1942 1810 1980
rect 1817 1942 1827 1980
rect 1829 1942 1866 1982
rect 1868 1980 1887 1982
rect 1868 1942 1876 1980
rect 1883 1942 1887 1980
rect 1931 1981 1951 1983
rect 1931 1943 1934 1981
rect 1941 1943 1951 1981
rect 1953 1943 1990 1983
rect 1992 1981 2011 1983
rect 1992 1943 2000 1981
rect 2007 1943 2011 1981
rect 2046 1981 2066 1983
rect 2046 1943 2049 1981
rect 2056 1943 2066 1981
rect 2068 1943 2105 1983
rect 2107 1981 2126 1983
rect 2107 1943 2115 1981
rect 2122 1943 2126 1981
rect 1084 1570 1104 1572
rect 1084 1532 1087 1570
rect 1094 1532 1104 1570
rect 1106 1532 1143 1572
rect 1145 1570 1164 1572
rect 1145 1532 1153 1570
rect 1160 1532 1164 1570
rect 1196 1508 1197 1528
rect 1199 1508 1200 1528
rect 1196 1304 1197 1324
rect 1199 1304 1200 1324
rect 1084 1262 1087 1300
rect 1094 1262 1104 1300
rect 1084 1260 1104 1262
rect 1106 1260 1143 1300
rect 1145 1262 1153 1300
rect 1160 1262 1164 1300
rect 1145 1260 1164 1262
rect 1084 1197 1104 1199
rect 1084 1159 1087 1197
rect 1094 1159 1104 1197
rect 1106 1159 1143 1199
rect 1145 1197 1164 1199
rect 1145 1159 1153 1197
rect 1160 1159 1164 1197
rect 1196 1135 1197 1155
rect 1199 1135 1200 1155
rect 1931 1687 1934 1725
rect 1941 1687 1951 1725
rect 1931 1685 1951 1687
rect 1953 1685 1990 1725
rect 1992 1687 2000 1725
rect 2007 1687 2011 1725
rect 1992 1685 2011 1687
rect 1547 1607 1567 1608
rect 1547 1604 1567 1605
rect 1570 1549 1610 1552
rect 1608 1542 1610 1549
rect 1570 1532 1610 1542
rect 1570 1493 1610 1530
rect 1570 1483 1610 1491
rect 1608 1476 1610 1483
rect 1570 1472 1610 1476
rect 1699 1437 1719 1438
rect 1547 1434 1567 1435
rect 1699 1434 1719 1435
rect 1547 1431 1567 1432
rect 1656 1379 1696 1382
rect 1551 1372 1571 1373
rect 1656 1372 1658 1379
rect 1551 1369 1571 1370
rect 1656 1362 1696 1372
rect 1656 1323 1696 1360
rect 1574 1314 1614 1317
rect 1612 1307 1614 1314
rect 1574 1297 1614 1307
rect 1656 1313 1696 1321
rect 1656 1306 1658 1313
rect 1656 1302 1696 1306
rect 1574 1258 1614 1295
rect 1699 1264 1719 1265
rect 1699 1261 1719 1262
rect 1574 1248 1614 1256
rect 1612 1241 1614 1248
rect 1574 1237 1614 1241
rect 2230 1805 2233 1843
rect 2240 1805 2250 1843
rect 2230 1803 2250 1805
rect 2252 1803 2289 1843
rect 2291 1805 2299 1843
rect 2306 1805 2310 1843
rect 2291 1803 2310 1805
rect 2230 1769 2250 1771
rect 2230 1731 2233 1769
rect 2240 1731 2250 1769
rect 2252 1731 2289 1771
rect 2291 1769 2310 1771
rect 2291 1731 2299 1769
rect 2306 1731 2310 1769
rect 2532 1770 2552 1772
rect 2532 1732 2535 1770
rect 2542 1732 2552 1770
rect 2554 1732 2591 1772
rect 2593 1770 2612 1772
rect 2593 1732 2601 1770
rect 2608 1732 2612 1770
rect 2360 1517 2361 1537
rect 2363 1517 2364 1537
rect 2230 1475 2233 1513
rect 2240 1475 2250 1513
rect 2230 1473 2250 1475
rect 2252 1473 2289 1513
rect 2291 1475 2299 1513
rect 2306 1475 2310 1513
rect 2291 1473 2310 1475
rect 2406 1476 2409 1514
rect 2416 1476 2426 1514
rect 2406 1474 2426 1476
rect 2428 1474 2465 1514
rect 2467 1476 2475 1514
rect 2482 1476 2486 1514
rect 2467 1474 2486 1476
rect 2230 1439 2250 1441
rect 2230 1401 2233 1439
rect 2240 1401 2250 1439
rect 2252 1401 2289 1441
rect 2291 1439 2310 1441
rect 2291 1401 2299 1439
rect 2306 1401 2310 1439
rect 2532 1476 2535 1514
rect 2542 1476 2552 1514
rect 2532 1474 2552 1476
rect 2554 1474 2591 1514
rect 2593 1476 2601 1514
rect 2608 1476 2612 1514
rect 2593 1474 2612 1476
rect 1551 1199 1571 1200
rect 1551 1196 1571 1197
rect 1690 1175 1710 1176
rect 1690 1172 1710 1173
rect 1647 1117 1687 1120
rect 1647 1110 1649 1117
rect 1647 1100 1687 1110
rect 1647 1061 1687 1098
rect 1647 1051 1687 1059
rect 1647 1044 1649 1051
rect 1647 1040 1687 1044
rect 1690 1002 1710 1003
rect 1690 999 1710 1000
rect 2230 1145 2233 1183
rect 2240 1145 2250 1183
rect 2230 1143 2250 1145
rect 2252 1143 2289 1183
rect 2291 1145 2299 1183
rect 2306 1145 2310 1183
rect 2291 1143 2310 1145
rect 2230 1109 2250 1111
rect 2230 1071 2233 1109
rect 2240 1071 2250 1109
rect 2252 1071 2289 1111
rect 2291 1109 2310 1111
rect 2291 1071 2299 1109
rect 2306 1071 2310 1109
rect 2532 1110 2552 1112
rect 2532 1072 2535 1110
rect 2542 1072 2552 1110
rect 2554 1072 2591 1112
rect 2593 1110 2612 1112
rect 2593 1072 2601 1110
rect 2608 1072 2612 1110
rect 2360 857 2361 877
rect 2363 857 2364 877
rect 2230 815 2233 853
rect 2240 815 2250 853
rect 2230 813 2250 815
rect 2252 813 2289 853
rect 2291 815 2299 853
rect 2306 815 2310 853
rect 2291 813 2310 815
rect 2406 816 2409 854
rect 2416 816 2426 854
rect 2406 814 2426 816
rect 2428 814 2465 854
rect 2467 816 2475 854
rect 2482 816 2486 854
rect 2467 814 2486 816
rect 2230 779 2250 781
rect 2230 741 2233 779
rect 2240 741 2250 779
rect 2252 741 2289 781
rect 2291 779 2310 781
rect 2291 741 2299 779
rect 2306 741 2310 779
rect 2532 816 2535 854
rect 2542 816 2552 854
rect 2532 814 2552 816
rect 2554 814 2591 854
rect 2593 816 2601 854
rect 2608 816 2612 854
rect 2593 814 2612 816
rect 185 126 225 129
rect 185 119 187 126
rect 185 109 225 119
rect 443 126 483 129
rect 185 70 225 107
rect 481 119 483 126
rect 443 109 483 119
rect 443 70 483 107
rect 185 60 225 68
rect 185 53 187 60
rect 185 49 225 53
rect 443 60 483 68
rect 481 53 483 60
rect 443 49 483 53
<< pdiffusion >>
rect 24 4259 64 4262
rect 24 4252 26 4259
rect 24 4242 64 4252
rect 272 4259 312 4262
rect 310 4252 312 4259
rect 272 4242 312 4252
rect 354 4259 394 4262
rect 354 4252 356 4259
rect 24 4225 64 4240
rect 24 4218 26 4225
rect 24 4203 64 4218
rect 272 4225 312 4240
rect 354 4242 394 4252
rect 602 4259 642 4262
rect 640 4252 642 4259
rect 602 4242 642 4252
rect 310 4218 312 4225
rect 272 4203 312 4218
rect 354 4225 394 4240
rect 354 4218 356 4225
rect 354 4203 394 4218
rect 602 4225 642 4240
rect 640 4218 642 4225
rect 602 4203 642 4218
rect 24 4192 64 4201
rect 24 4185 26 4192
rect 24 4182 64 4185
rect 272 4192 312 4201
rect 310 4185 312 4192
rect 272 4182 312 4185
rect 354 4192 394 4201
rect 354 4185 356 4192
rect 354 4182 394 4185
rect 602 4192 642 4201
rect 640 4185 642 4192
rect 602 4182 642 4185
rect 270 4131 320 4132
rect 270 4128 320 4129
rect 273 4083 313 4086
rect 311 4076 313 4083
rect 273 4066 313 4076
rect 273 4049 313 4064
rect 311 4042 313 4049
rect 273 4027 313 4042
rect 273 4016 313 4025
rect 311 4009 313 4016
rect 273 4006 313 4009
rect 273 3957 313 3960
rect 311 3950 313 3957
rect 273 3940 313 3950
rect 355 3957 395 3960
rect 355 3950 357 3957
rect 273 3923 313 3938
rect 355 3940 395 3950
rect 311 3916 313 3923
rect 273 3901 313 3916
rect 355 3923 395 3938
rect 355 3916 357 3923
rect 355 3901 395 3916
rect 273 3890 313 3899
rect 311 3883 313 3890
rect 273 3880 313 3883
rect 355 3890 395 3899
rect 355 3883 357 3890
rect 355 3880 395 3883
rect 2230 3909 2250 3911
rect 2230 3871 2233 3909
rect 2240 3871 2250 3909
rect 2252 3909 2289 3911
rect 2252 3871 2267 3909
rect 2274 3871 2289 3909
rect 2291 3909 2310 3911
rect 2291 3871 2300 3909
rect 2307 3871 2310 3909
rect 1182 3623 1232 3624
rect 1182 3620 1232 3621
rect 1185 3565 1225 3568
rect 1223 3558 1225 3565
rect 1185 3548 1225 3558
rect 1185 3531 1225 3546
rect 1223 3524 1225 3531
rect 1185 3509 1225 3524
rect 24 3302 64 3305
rect 24 3295 26 3302
rect 24 3285 64 3295
rect 272 3302 312 3305
rect 310 3295 312 3302
rect 272 3285 312 3295
rect 354 3302 394 3305
rect 354 3295 356 3302
rect 24 3268 64 3283
rect 24 3261 26 3268
rect 24 3246 64 3261
rect 272 3268 312 3283
rect 354 3285 394 3295
rect 602 3302 642 3305
rect 640 3295 642 3302
rect 602 3285 642 3295
rect 310 3261 312 3268
rect 272 3246 312 3261
rect 354 3268 394 3283
rect 354 3261 356 3268
rect 354 3246 394 3261
rect 602 3268 642 3283
rect 1185 3498 1225 3507
rect 1223 3491 1225 3498
rect 1185 3488 1225 3491
rect 1182 3450 1232 3451
rect 1182 3447 1232 3448
rect 1931 3460 1934 3498
rect 1941 3460 1951 3498
rect 1931 3458 1951 3460
rect 1953 3460 1968 3498
rect 1975 3460 1990 3498
rect 1953 3458 1990 3460
rect 1992 3460 2001 3498
rect 2008 3460 2011 3498
rect 1992 3458 2011 3460
rect 1807 3415 1827 3417
rect 1185 3400 1225 3403
rect 1223 3393 1225 3400
rect 1185 3383 1225 3393
rect 1185 3366 1225 3381
rect 1223 3359 1225 3366
rect 1185 3344 1225 3359
rect 1807 3377 1810 3415
rect 1817 3377 1827 3415
rect 1829 3415 1866 3417
rect 1829 3377 1844 3415
rect 1851 3377 1866 3415
rect 1868 3415 1887 3417
rect 1868 3377 1877 3415
rect 1884 3377 1887 3415
rect 1185 3333 1225 3342
rect 1223 3326 1225 3333
rect 1185 3323 1225 3326
rect 1183 3290 1233 3291
rect 1183 3287 1233 3288
rect 640 3261 642 3268
rect 602 3246 642 3261
rect 24 3235 64 3244
rect 24 3228 26 3235
rect 24 3225 64 3228
rect 272 3235 312 3244
rect 310 3228 312 3235
rect 272 3225 312 3228
rect 354 3235 394 3244
rect 354 3228 356 3235
rect 354 3225 394 3228
rect 602 3235 642 3244
rect 640 3228 642 3235
rect 602 3225 642 3228
rect 270 3174 320 3175
rect 270 3171 320 3172
rect 273 3126 313 3129
rect 311 3119 313 3126
rect 273 3109 313 3119
rect 273 3092 313 3107
rect 311 3085 313 3092
rect 273 3070 313 3085
rect 273 3059 313 3068
rect 311 3052 313 3059
rect 273 3049 313 3052
rect 1931 3414 1951 3416
rect 1931 3376 1934 3414
rect 1941 3376 1951 3414
rect 1953 3414 1990 3416
rect 1953 3376 1968 3414
rect 1975 3376 1990 3414
rect 1992 3414 2011 3416
rect 1992 3376 2001 3414
rect 2008 3376 2011 3414
rect 2046 3414 2066 3416
rect 2046 3376 2049 3414
rect 2056 3376 2066 3414
rect 2068 3414 2105 3416
rect 2068 3376 2083 3414
rect 2090 3376 2105 3414
rect 2107 3414 2126 3416
rect 2107 3376 2116 3414
rect 2123 3376 2126 3414
rect 2230 3625 2233 3663
rect 2240 3625 2250 3663
rect 2230 3623 2250 3625
rect 2252 3625 2267 3663
rect 2274 3625 2289 3663
rect 2252 3623 2289 3625
rect 2291 3625 2300 3663
rect 2307 3625 2310 3663
rect 2291 3623 2310 3625
rect 2532 3626 2535 3664
rect 2542 3626 2552 3664
rect 2532 3624 2552 3626
rect 2554 3626 2569 3664
rect 2576 3626 2591 3664
rect 2554 3624 2591 3626
rect 2593 3626 2602 3664
rect 2609 3626 2612 3664
rect 2593 3624 2612 3626
rect 2230 3579 2250 3581
rect 2230 3541 2233 3579
rect 2240 3541 2250 3579
rect 2252 3579 2289 3581
rect 2252 3541 2267 3579
rect 2274 3541 2289 3579
rect 2291 3579 2310 3581
rect 2291 3541 2300 3579
rect 2307 3541 2310 3579
rect 2360 3539 2361 3589
rect 2363 3539 2364 3589
rect 2406 3580 2426 3582
rect 2406 3542 2409 3580
rect 2416 3542 2426 3580
rect 2428 3580 2465 3582
rect 2428 3542 2443 3580
rect 2450 3542 2465 3580
rect 2467 3580 2486 3582
rect 2467 3542 2476 3580
rect 2483 3542 2486 3580
rect 2532 3580 2552 3582
rect 2532 3542 2535 3580
rect 2542 3542 2552 3580
rect 2554 3580 2591 3582
rect 2554 3542 2569 3580
rect 2576 3542 2591 3580
rect 2593 3580 2612 3582
rect 2593 3542 2602 3580
rect 2609 3542 2612 3580
rect 2230 3295 2233 3333
rect 2240 3295 2250 3333
rect 2230 3293 2250 3295
rect 2252 3295 2267 3333
rect 2274 3295 2289 3333
rect 2252 3293 2289 3295
rect 2291 3295 2300 3333
rect 2307 3295 2310 3333
rect 2291 3293 2310 3295
rect 2230 3249 2250 3251
rect 2230 3211 2233 3249
rect 2240 3211 2250 3249
rect 2252 3249 2289 3251
rect 2252 3211 2267 3249
rect 2274 3211 2289 3249
rect 2291 3249 2310 3251
rect 2291 3211 2300 3249
rect 2307 3211 2310 3249
rect 737 3102 740 3140
rect 747 3102 757 3140
rect 737 3100 757 3102
rect 759 3102 774 3140
rect 781 3102 796 3140
rect 759 3100 796 3102
rect 798 3102 807 3140
rect 814 3102 817 3140
rect 798 3100 817 3102
rect 1194 3179 1234 3182
rect 1232 3172 1234 3179
rect 1194 3162 1234 3172
rect 861 3103 864 3141
rect 871 3103 881 3141
rect 861 3101 881 3103
rect 883 3103 898 3141
rect 905 3103 920 3141
rect 883 3101 920 3103
rect 922 3103 931 3141
rect 938 3103 941 3141
rect 922 3101 941 3103
rect 976 3103 979 3141
rect 986 3103 996 3141
rect 976 3101 996 3103
rect 998 3103 1013 3141
rect 1020 3103 1035 3141
rect 998 3101 1035 3103
rect 1037 3103 1046 3141
rect 1053 3103 1056 3141
rect 1037 3101 1056 3103
rect 1194 3145 1234 3160
rect 1232 3138 1234 3145
rect 1194 3123 1234 3138
rect 861 3057 881 3059
rect 861 3019 864 3057
rect 871 3019 881 3057
rect 883 3057 920 3059
rect 883 3019 898 3057
rect 905 3019 920 3057
rect 922 3057 941 3059
rect 922 3019 931 3057
rect 938 3019 941 3057
rect 273 3000 313 3003
rect 311 2993 313 3000
rect 273 2983 313 2993
rect 355 3000 395 3003
rect 355 2993 357 3000
rect 273 2966 313 2981
rect 355 2983 395 2993
rect 311 2959 313 2966
rect 273 2944 313 2959
rect 355 2966 395 2981
rect 355 2959 357 2966
rect 355 2944 395 2959
rect 273 2933 313 2942
rect 311 2926 313 2933
rect 273 2923 313 2926
rect 355 2933 395 2942
rect 355 2926 357 2933
rect 355 2923 395 2926
rect 24 2823 64 2826
rect 24 2816 26 2823
rect 24 2806 64 2816
rect 272 2823 312 2826
rect 310 2816 312 2823
rect 272 2806 312 2816
rect 354 2823 394 2826
rect 354 2816 356 2823
rect 24 2789 64 2804
rect 24 2782 26 2789
rect 24 2767 64 2782
rect 272 2789 312 2804
rect 354 2806 394 2816
rect 602 2823 642 2826
rect 640 2816 642 2823
rect 602 2806 642 2816
rect 310 2782 312 2789
rect 272 2767 312 2782
rect 354 2789 394 2804
rect 354 2782 356 2789
rect 354 2767 394 2782
rect 602 2789 642 2804
rect 640 2782 642 2789
rect 602 2767 642 2782
rect 24 2756 64 2765
rect 24 2749 26 2756
rect 24 2746 64 2749
rect 272 2756 312 2765
rect 310 2749 312 2756
rect 272 2746 312 2749
rect 354 2756 394 2765
rect 354 2749 356 2756
rect 354 2746 394 2749
rect 602 2756 642 2765
rect 640 2749 642 2756
rect 602 2746 642 2749
rect 270 2695 320 2696
rect 270 2692 320 2693
rect 273 2647 313 2650
rect 311 2640 313 2647
rect 273 2630 313 2640
rect 273 2613 313 2628
rect 311 2606 313 2613
rect 273 2591 313 2606
rect 273 2580 313 2589
rect 311 2573 313 2580
rect 273 2570 313 2573
rect 723 2884 763 2887
rect 723 2877 725 2884
rect 723 2867 763 2877
rect 723 2850 763 2865
rect 723 2843 725 2850
rect 723 2828 763 2843
rect 723 2817 763 2826
rect 723 2810 725 2817
rect 723 2807 763 2810
rect 715 2774 765 2775
rect 715 2771 765 2772
rect 1194 3112 1234 3121
rect 1232 3105 1234 3112
rect 1194 3102 1234 3105
rect 1192 3069 1242 3070
rect 1192 3066 1242 3067
rect 1807 2982 1810 3020
rect 1817 2982 1827 3020
rect 1807 2980 1827 2982
rect 1829 2982 1844 3020
rect 1851 2982 1866 3020
rect 1829 2980 1866 2982
rect 1868 2982 1877 3020
rect 1884 2982 1887 3020
rect 1868 2980 1887 2982
rect 1195 2974 1235 2977
rect 1233 2967 1235 2974
rect 1195 2957 1235 2967
rect 1195 2940 1235 2955
rect 1233 2933 1235 2940
rect 1195 2918 1235 2933
rect 1195 2907 1235 2916
rect 1233 2900 1235 2907
rect 1195 2897 1235 2900
rect 1931 2983 1934 3021
rect 1941 2983 1951 3021
rect 1931 2981 1951 2983
rect 1953 2983 1968 3021
rect 1975 2983 1990 3021
rect 1953 2981 1990 2983
rect 1992 2983 2001 3021
rect 2008 2983 2011 3021
rect 1992 2981 2011 2983
rect 2046 2983 2049 3021
rect 2056 2983 2066 3021
rect 2046 2981 2066 2983
rect 2068 2983 2083 3021
rect 2090 2983 2105 3021
rect 2068 2981 2105 2983
rect 2107 2983 2116 3021
rect 2123 2983 2126 3021
rect 2107 2981 2126 2983
rect 1931 2937 1951 2939
rect 1931 2899 1934 2937
rect 1941 2899 1951 2937
rect 1953 2937 1990 2939
rect 1953 2899 1968 2937
rect 1975 2899 1990 2937
rect 1992 2937 2011 2939
rect 1992 2899 2001 2937
rect 2008 2899 2011 2937
rect 1193 2864 1243 2865
rect 1193 2861 1243 2862
rect 1193 2783 1243 2784
rect 1193 2780 1243 2781
rect 273 2521 313 2524
rect 311 2514 313 2521
rect 273 2504 313 2514
rect 355 2521 395 2524
rect 355 2514 357 2521
rect 273 2487 313 2502
rect 355 2504 395 2514
rect 311 2480 313 2487
rect 273 2465 313 2480
rect 355 2487 395 2502
rect 355 2480 357 2487
rect 355 2465 395 2480
rect 273 2454 313 2463
rect 311 2447 313 2454
rect 273 2444 313 2447
rect 355 2454 395 2463
rect 355 2447 357 2454
rect 355 2444 395 2447
rect 24 2344 64 2347
rect 24 2337 26 2344
rect 24 2327 64 2337
rect 272 2344 312 2347
rect 310 2337 312 2344
rect 272 2327 312 2337
rect 354 2344 394 2347
rect 354 2337 356 2344
rect 24 2310 64 2325
rect 24 2303 26 2310
rect 24 2288 64 2303
rect 272 2310 312 2325
rect 354 2327 394 2337
rect 602 2344 642 2347
rect 640 2337 642 2344
rect 602 2327 642 2337
rect 310 2303 312 2310
rect 272 2288 312 2303
rect 354 2310 394 2325
rect 354 2303 356 2310
rect 354 2288 394 2303
rect 602 2310 642 2325
rect 640 2303 642 2310
rect 602 2288 642 2303
rect 24 2277 64 2286
rect 24 2270 26 2277
rect 24 2267 64 2270
rect 272 2277 312 2286
rect 310 2270 312 2277
rect 272 2267 312 2270
rect 354 2277 394 2286
rect 354 2270 356 2277
rect 354 2267 394 2270
rect 602 2277 642 2286
rect 640 2270 642 2277
rect 602 2267 642 2270
rect 270 2216 320 2217
rect 270 2213 320 2214
rect 273 2168 313 2171
rect 311 2161 313 2168
rect 273 2151 313 2161
rect 273 2134 313 2149
rect 311 2127 313 2134
rect 273 2112 313 2127
rect 273 2101 313 2110
rect 311 2094 313 2101
rect 273 2091 313 2094
rect 1196 2725 1236 2728
rect 1234 2718 1236 2725
rect 1196 2708 1236 2718
rect 1196 2691 1236 2706
rect 1234 2684 1236 2691
rect 1196 2669 1236 2684
rect 715 2645 765 2646
rect 715 2642 765 2643
rect 1196 2658 1236 2667
rect 1234 2651 1236 2658
rect 1196 2648 1236 2651
rect 1193 2610 1243 2611
rect 723 2607 763 2610
rect 723 2600 725 2607
rect 723 2591 763 2600
rect 1193 2607 1243 2608
rect 723 2574 763 2589
rect 723 2567 725 2574
rect 723 2552 763 2567
rect 723 2540 763 2550
rect 723 2533 725 2540
rect 723 2530 763 2533
rect 737 2315 757 2317
rect 737 2277 740 2315
rect 747 2277 757 2315
rect 759 2315 796 2317
rect 759 2277 774 2315
rect 781 2277 796 2315
rect 798 2315 817 2317
rect 798 2277 807 2315
rect 814 2277 817 2315
rect 861 2360 864 2398
rect 871 2360 881 2398
rect 861 2358 881 2360
rect 883 2360 898 2398
rect 905 2360 920 2398
rect 883 2358 920 2360
rect 922 2360 931 2398
rect 938 2360 941 2398
rect 922 2358 941 2360
rect 861 2314 881 2316
rect 861 2276 864 2314
rect 871 2276 881 2314
rect 883 2314 920 2316
rect 883 2276 898 2314
rect 905 2276 920 2314
rect 922 2314 941 2316
rect 922 2276 931 2314
rect 938 2276 941 2314
rect 976 2314 996 2316
rect 976 2276 979 2314
rect 986 2276 996 2314
rect 998 2314 1035 2316
rect 998 2276 1013 2314
rect 1020 2276 1035 2314
rect 1037 2314 1056 2316
rect 1037 2276 1046 2314
rect 1053 2276 1056 2314
rect 1091 2314 1111 2316
rect 1091 2276 1094 2314
rect 1101 2276 1111 2314
rect 1113 2314 1150 2316
rect 1113 2276 1128 2314
rect 1135 2276 1150 2314
rect 1152 2314 1171 2316
rect 1152 2276 1161 2314
rect 1168 2276 1171 2314
rect 273 2042 313 2045
rect 311 2035 313 2042
rect 273 2025 313 2035
rect 355 2042 395 2045
rect 355 2035 357 2042
rect 273 2008 313 2023
rect 355 2025 395 2035
rect 311 2001 313 2008
rect 273 1986 313 2001
rect 355 2008 395 2023
rect 355 2001 357 2008
rect 355 1986 395 2001
rect 273 1975 313 1984
rect 311 1968 313 1975
rect 273 1965 313 1968
rect 355 1975 395 1984
rect 355 1968 357 1975
rect 355 1965 395 1968
rect 24 1865 64 1868
rect 24 1858 26 1865
rect 24 1848 64 1858
rect 272 1865 312 1868
rect 310 1858 312 1865
rect 272 1848 312 1858
rect 354 1865 394 1868
rect 354 1858 356 1865
rect 24 1831 64 1846
rect 24 1824 26 1831
rect 24 1809 64 1824
rect 272 1831 312 1846
rect 354 1848 394 1858
rect 602 1865 642 1868
rect 640 1858 642 1865
rect 602 1848 642 1858
rect 310 1824 312 1831
rect 272 1809 312 1824
rect 354 1831 394 1846
rect 354 1824 356 1831
rect 354 1809 394 1824
rect 602 1831 642 1846
rect 640 1824 642 1831
rect 602 1809 642 1824
rect 24 1798 64 1807
rect 24 1791 26 1798
rect 24 1788 64 1791
rect 272 1798 312 1807
rect 310 1791 312 1798
rect 272 1788 312 1791
rect 354 1798 394 1807
rect 354 1791 356 1798
rect 354 1788 394 1791
rect 602 1798 642 1807
rect 1203 2274 1204 2324
rect 1206 2274 1207 2324
rect 1315 2733 1365 2734
rect 1315 2730 1365 2731
rect 2230 2965 2233 3003
rect 2240 2965 2250 3003
rect 2230 2963 2250 2965
rect 2252 2965 2267 3003
rect 2274 2965 2289 3003
rect 2252 2963 2289 2965
rect 2291 2965 2300 3003
rect 2307 2965 2310 3003
rect 2291 2963 2310 2965
rect 2532 2966 2535 3004
rect 2542 2966 2552 3004
rect 2532 2964 2552 2966
rect 2554 2966 2569 3004
rect 2576 2966 2591 3004
rect 2554 2964 2591 2966
rect 2593 2966 2602 3004
rect 2609 2966 2612 3004
rect 2593 2964 2612 2966
rect 2230 2919 2250 2921
rect 2230 2881 2233 2919
rect 2240 2881 2250 2919
rect 2252 2919 2289 2921
rect 2252 2881 2267 2919
rect 2274 2881 2289 2919
rect 2291 2919 2310 2921
rect 2291 2881 2300 2919
rect 2307 2881 2310 2919
rect 2360 2879 2361 2929
rect 2363 2879 2364 2929
rect 2406 2920 2426 2922
rect 2406 2882 2409 2920
rect 2416 2882 2426 2920
rect 2428 2920 2465 2922
rect 2428 2882 2443 2920
rect 2450 2882 2465 2920
rect 2467 2920 2486 2922
rect 2467 2882 2476 2920
rect 2483 2882 2486 2920
rect 2532 2920 2552 2922
rect 2532 2882 2535 2920
rect 2542 2882 2552 2920
rect 2554 2920 2591 2922
rect 2554 2882 2569 2920
rect 2576 2882 2591 2920
rect 2593 2920 2612 2922
rect 2593 2882 2602 2920
rect 2609 2882 2612 2920
rect 1322 2675 1362 2678
rect 1322 2668 1324 2675
rect 1322 2658 1362 2668
rect 1322 2641 1362 2656
rect 1322 2634 1324 2641
rect 1322 2619 1362 2634
rect 2230 2635 2233 2673
rect 2240 2635 2250 2673
rect 2230 2633 2250 2635
rect 2252 2635 2267 2673
rect 2274 2635 2289 2673
rect 2252 2633 2289 2635
rect 2291 2635 2300 2673
rect 2307 2635 2310 2673
rect 2291 2633 2310 2635
rect 1322 2608 1362 2617
rect 1322 2601 1324 2608
rect 1322 2598 1362 2601
rect 1315 2560 1365 2561
rect 1315 2557 1365 2558
rect 640 1791 642 1798
rect 602 1788 642 1791
rect 270 1737 320 1738
rect 270 1734 320 1735
rect 273 1689 313 1692
rect 311 1682 313 1689
rect 273 1672 313 1682
rect 273 1655 313 1670
rect 311 1648 313 1655
rect 273 1633 313 1648
rect 273 1622 313 1631
rect 311 1615 313 1622
rect 273 1612 313 1615
rect 737 1976 740 2014
rect 747 1976 757 2014
rect 737 1974 757 1976
rect 759 1976 774 2014
rect 781 1976 796 2014
rect 759 1974 796 1976
rect 798 1976 807 2014
rect 814 1976 817 2014
rect 798 1974 817 1976
rect 861 1977 864 2015
rect 871 1977 881 2015
rect 861 1975 881 1977
rect 883 1977 898 2015
rect 905 1977 920 2015
rect 883 1975 920 1977
rect 922 1977 931 2015
rect 938 1977 941 2015
rect 922 1975 941 1977
rect 976 1977 979 2015
rect 986 1977 996 2015
rect 976 1975 996 1977
rect 998 1977 1013 2015
rect 1020 1977 1035 2015
rect 998 1975 1035 1977
rect 1037 1977 1046 2015
rect 1053 1977 1056 2015
rect 1037 1975 1056 1977
rect 861 1931 881 1933
rect 861 1893 864 1931
rect 871 1893 881 1931
rect 883 1931 920 1933
rect 883 1893 898 1931
rect 905 1893 920 1931
rect 922 1931 941 1933
rect 922 1893 931 1931
rect 938 1893 941 1931
rect 273 1563 313 1566
rect 311 1556 313 1563
rect 273 1546 313 1556
rect 355 1563 395 1566
rect 355 1556 357 1563
rect 273 1529 313 1544
rect 355 1546 395 1556
rect 311 1522 313 1529
rect 273 1507 313 1522
rect 355 1529 395 1544
rect 355 1522 357 1529
rect 355 1507 395 1522
rect 273 1496 313 1505
rect 311 1489 313 1496
rect 273 1486 313 1489
rect 355 1496 395 1505
rect 355 1489 357 1496
rect 355 1486 395 1489
rect 24 1386 64 1389
rect 24 1379 26 1386
rect 24 1369 64 1379
rect 272 1386 312 1389
rect 310 1379 312 1386
rect 272 1369 312 1379
rect 354 1386 394 1389
rect 354 1379 356 1386
rect 24 1352 64 1367
rect 24 1345 26 1352
rect 24 1330 64 1345
rect 272 1352 312 1367
rect 354 1369 394 1379
rect 602 1386 642 1389
rect 640 1379 642 1386
rect 602 1369 642 1379
rect 310 1345 312 1352
rect 272 1330 312 1345
rect 354 1352 394 1367
rect 354 1345 356 1352
rect 354 1330 394 1345
rect 602 1352 642 1367
rect 640 1345 642 1352
rect 602 1330 642 1345
rect 24 1319 64 1328
rect 24 1312 26 1319
rect 24 1309 64 1312
rect 272 1319 312 1328
rect 310 1312 312 1319
rect 272 1309 312 1312
rect 354 1319 394 1328
rect 354 1312 356 1319
rect 354 1309 394 1312
rect 602 1319 642 1328
rect 640 1312 642 1319
rect 602 1309 642 1312
rect 270 1258 320 1259
rect 270 1255 320 1256
rect 273 1210 313 1213
rect 311 1203 313 1210
rect 273 1193 313 1203
rect 273 1176 313 1191
rect 311 1169 313 1176
rect 273 1154 313 1169
rect 273 1143 313 1152
rect 311 1136 313 1143
rect 273 1133 313 1136
rect 723 1758 763 1761
rect 723 1751 725 1758
rect 723 1741 763 1751
rect 723 1724 763 1739
rect 723 1717 725 1724
rect 723 1702 763 1717
rect 723 1691 763 1700
rect 723 1684 725 1691
rect 723 1681 763 1684
rect 715 1648 765 1649
rect 715 1645 765 1646
rect 273 1084 313 1087
rect 311 1077 313 1084
rect 273 1067 313 1077
rect 355 1084 395 1087
rect 355 1077 357 1084
rect 273 1050 313 1065
rect 355 1067 395 1077
rect 311 1043 313 1050
rect 273 1028 313 1043
rect 355 1050 395 1065
rect 355 1043 357 1050
rect 355 1028 395 1043
rect 273 1017 313 1026
rect 311 1010 313 1017
rect 273 1007 313 1010
rect 355 1017 395 1026
rect 355 1010 357 1017
rect 355 1007 395 1010
rect 24 907 64 910
rect 24 900 26 907
rect 24 890 64 900
rect 272 907 312 910
rect 310 900 312 907
rect 272 890 312 900
rect 354 907 394 910
rect 354 900 356 907
rect 24 873 64 888
rect 24 866 26 873
rect 24 851 64 866
rect 272 873 312 888
rect 354 890 394 900
rect 602 907 642 910
rect 640 900 642 907
rect 602 890 642 900
rect 310 866 312 873
rect 272 851 312 866
rect 354 873 394 888
rect 354 866 356 873
rect 354 851 394 866
rect 602 873 642 888
rect 640 866 642 873
rect 602 851 642 866
rect 24 840 64 849
rect 24 833 26 840
rect 24 830 64 833
rect 272 840 312 849
rect 310 833 312 840
rect 272 830 312 833
rect 354 840 394 849
rect 354 833 356 840
rect 354 830 394 833
rect 602 840 642 849
rect 640 833 642 840
rect 602 830 642 833
rect 270 779 320 780
rect 270 776 320 777
rect 273 731 313 734
rect 311 724 313 731
rect 273 714 313 724
rect 273 697 313 712
rect 311 690 313 697
rect 273 675 313 690
rect 273 664 313 673
rect 311 657 313 664
rect 273 654 313 657
rect 273 605 313 608
rect 311 598 313 605
rect 273 588 313 598
rect 355 605 395 608
rect 355 598 357 605
rect 273 571 313 586
rect 355 588 395 598
rect 311 564 313 571
rect 273 549 313 564
rect 355 571 395 586
rect 355 564 357 571
rect 355 549 395 564
rect 273 538 313 547
rect 311 531 313 538
rect 273 528 313 531
rect 355 538 395 547
rect 355 531 357 538
rect 355 528 395 531
rect 24 428 64 431
rect 24 421 26 428
rect 24 411 64 421
rect 272 428 312 431
rect 310 421 312 428
rect 272 411 312 421
rect 354 428 394 431
rect 354 421 356 428
rect 24 394 64 409
rect 24 387 26 394
rect 24 372 64 387
rect 272 394 312 409
rect 354 411 394 421
rect 602 428 642 431
rect 640 421 642 428
rect 602 411 642 421
rect 310 387 312 394
rect 272 372 312 387
rect 354 394 394 409
rect 354 387 356 394
rect 354 372 394 387
rect 602 394 642 409
rect 640 387 642 394
rect 602 372 642 387
rect 24 361 64 370
rect 24 354 26 361
rect 24 351 64 354
rect 272 361 312 370
rect 310 354 312 361
rect 272 351 312 354
rect 354 361 394 370
rect 354 354 356 361
rect 354 351 394 354
rect 602 361 642 370
rect 640 354 642 361
rect 602 351 642 354
rect 270 300 320 301
rect 270 297 320 298
rect 273 252 313 255
rect 311 245 313 252
rect 273 235 313 245
rect 273 218 313 233
rect 311 211 313 218
rect 273 196 313 211
rect 273 185 313 194
rect 311 178 313 185
rect 273 175 313 178
rect 1091 2030 1094 2068
rect 1101 2030 1111 2068
rect 1091 2028 1111 2030
rect 1113 2030 1128 2068
rect 1135 2030 1150 2068
rect 1113 2028 1150 2030
rect 1152 2030 1161 2068
rect 1168 2030 1171 2068
rect 1152 2028 1171 2030
rect 1203 2020 1204 2070
rect 1206 2020 1207 2070
rect 2230 2589 2250 2591
rect 2230 2551 2233 2589
rect 2240 2551 2250 2589
rect 2252 2589 2289 2591
rect 2252 2551 2267 2589
rect 2274 2551 2289 2589
rect 2291 2589 2310 2591
rect 2291 2551 2300 2589
rect 2307 2551 2310 2589
rect 1378 2378 1428 2379
rect 1378 2375 1428 2376
rect 1385 2320 1425 2323
rect 1385 2313 1387 2320
rect 1385 2303 1425 2313
rect 1931 2334 1934 2372
rect 1941 2334 1951 2372
rect 1931 2332 1951 2334
rect 1953 2334 1968 2372
rect 1975 2334 1990 2372
rect 1953 2332 1990 2334
rect 1992 2334 2001 2372
rect 2008 2334 2011 2372
rect 1992 2332 2011 2334
rect 1385 2286 1425 2301
rect 1385 2279 1387 2286
rect 1385 2264 1425 2279
rect 1807 2289 1827 2291
rect 1385 2253 1425 2262
rect 1385 2246 1387 2253
rect 1385 2243 1425 2246
rect 1807 2251 1810 2289
rect 1817 2251 1827 2289
rect 1829 2289 1866 2291
rect 1829 2251 1844 2289
rect 1851 2251 1866 2289
rect 1868 2289 1887 2291
rect 1868 2251 1877 2289
rect 1884 2251 1887 2289
rect 1378 2205 1428 2206
rect 1644 2208 1694 2209
rect 1378 2202 1428 2203
rect 1644 2205 1694 2206
rect 1931 2288 1951 2290
rect 1931 2250 1934 2288
rect 1941 2250 1951 2288
rect 1953 2288 1990 2290
rect 1953 2250 1968 2288
rect 1975 2250 1990 2288
rect 1992 2288 2011 2290
rect 1992 2250 2001 2288
rect 2008 2250 2011 2288
rect 1382 2143 1432 2144
rect 1647 2150 1687 2153
rect 1685 2143 1687 2150
rect 1382 2140 1432 2141
rect 1647 2133 1687 2143
rect 1647 2116 1687 2131
rect 1685 2109 1687 2116
rect 1647 2094 1687 2109
rect 1389 2085 1429 2088
rect 1389 2078 1391 2085
rect 1389 2068 1429 2078
rect 1389 2051 1429 2066
rect 1389 2044 1391 2051
rect 1389 2029 1429 2044
rect 1647 2083 1687 2092
rect 1685 2076 1687 2083
rect 1647 2073 1687 2076
rect 2046 2288 2066 2290
rect 2046 2250 2049 2288
rect 2056 2250 2066 2288
rect 2068 2288 2105 2290
rect 2068 2250 2083 2288
rect 2090 2250 2105 2288
rect 2107 2288 2126 2290
rect 2107 2250 2116 2288
rect 2123 2250 2126 2288
rect 1644 2035 1694 2036
rect 1389 2018 1429 2027
rect 1389 2011 1391 2018
rect 1389 2008 1429 2011
rect 1644 2032 1694 2033
rect 1091 1968 1111 1970
rect 1091 1930 1094 1968
rect 1101 1930 1111 1968
rect 1113 1968 1150 1970
rect 1113 1930 1128 1968
rect 1135 1930 1150 1968
rect 1152 1968 1171 1970
rect 1152 1930 1161 1968
rect 1168 1930 1171 1968
rect 1203 1928 1204 1978
rect 1206 1928 1207 1978
rect 2230 2305 2233 2343
rect 2240 2305 2250 2343
rect 2230 2303 2250 2305
rect 2252 2305 2267 2343
rect 2274 2305 2289 2343
rect 2252 2303 2289 2305
rect 2291 2305 2300 2343
rect 2307 2305 2310 2343
rect 2291 2303 2310 2305
rect 2532 2306 2535 2344
rect 2542 2306 2552 2344
rect 2532 2304 2552 2306
rect 2554 2306 2569 2344
rect 2576 2306 2591 2344
rect 2554 2304 2591 2306
rect 2593 2306 2602 2344
rect 2609 2306 2612 2344
rect 2593 2304 2612 2306
rect 2230 2259 2250 2261
rect 2230 2221 2233 2259
rect 2240 2221 2250 2259
rect 2252 2259 2289 2261
rect 2252 2221 2267 2259
rect 2274 2221 2289 2259
rect 2291 2259 2310 2261
rect 2291 2221 2300 2259
rect 2307 2221 2310 2259
rect 2360 2219 2361 2269
rect 2363 2219 2364 2269
rect 2406 2260 2426 2262
rect 2406 2222 2409 2260
rect 2416 2222 2426 2260
rect 2428 2260 2465 2262
rect 2428 2222 2443 2260
rect 2450 2222 2465 2260
rect 2467 2260 2486 2262
rect 2467 2222 2476 2260
rect 2483 2222 2486 2260
rect 2532 2260 2552 2262
rect 2532 2222 2535 2260
rect 2542 2222 2552 2260
rect 2554 2260 2591 2262
rect 2554 2222 2569 2260
rect 2576 2222 2591 2260
rect 2593 2260 2612 2262
rect 2593 2222 2602 2260
rect 2609 2222 2612 2260
rect 1382 1970 1432 1971
rect 1382 1967 1432 1968
rect 1088 1647 1091 1685
rect 1098 1647 1108 1685
rect 1088 1645 1108 1647
rect 1110 1647 1125 1685
rect 1132 1647 1147 1685
rect 1110 1645 1147 1647
rect 1149 1647 1158 1685
rect 1165 1647 1168 1685
rect 1149 1645 1168 1647
rect 1200 1637 1201 1687
rect 1203 1637 1204 1687
rect 2230 1975 2233 2013
rect 2240 1975 2250 2013
rect 2230 1973 2250 1975
rect 2252 1975 2267 2013
rect 2274 1975 2289 2013
rect 2252 1973 2289 1975
rect 2291 1975 2300 2013
rect 2307 1975 2310 2013
rect 2291 1973 2310 1975
rect 1084 1446 1087 1484
rect 1094 1446 1104 1484
rect 1084 1444 1104 1446
rect 1106 1446 1121 1484
rect 1128 1446 1143 1484
rect 1106 1444 1143 1446
rect 1145 1446 1154 1484
rect 1161 1446 1164 1484
rect 1145 1444 1164 1446
rect 1196 1436 1197 1486
rect 1199 1436 1200 1486
rect 1084 1386 1104 1388
rect 1084 1348 1087 1386
rect 1094 1348 1104 1386
rect 1106 1386 1143 1388
rect 1106 1348 1121 1386
rect 1128 1348 1143 1386
rect 1145 1386 1164 1388
rect 1145 1348 1154 1386
rect 1161 1348 1164 1386
rect 1196 1346 1197 1396
rect 1199 1346 1200 1396
rect 1084 1073 1087 1111
rect 1094 1073 1104 1111
rect 1084 1071 1104 1073
rect 1106 1073 1121 1111
rect 1128 1073 1143 1111
rect 1106 1071 1143 1073
rect 1145 1073 1154 1111
rect 1161 1073 1164 1111
rect 1145 1071 1164 1073
rect 1196 1063 1197 1113
rect 1199 1063 1200 1113
rect 1807 1856 1810 1894
rect 1817 1856 1827 1894
rect 1807 1854 1827 1856
rect 1829 1856 1844 1894
rect 1851 1856 1866 1894
rect 1829 1854 1866 1856
rect 1868 1856 1877 1894
rect 1884 1856 1887 1894
rect 1868 1854 1887 1856
rect 2230 1929 2250 1931
rect 1931 1857 1934 1895
rect 1941 1857 1951 1895
rect 1931 1855 1951 1857
rect 1953 1857 1968 1895
rect 1975 1857 1990 1895
rect 1953 1855 1990 1857
rect 1992 1857 2001 1895
rect 2008 1857 2011 1895
rect 1992 1855 2011 1857
rect 2046 1857 2049 1895
rect 2056 1857 2066 1895
rect 2046 1855 2066 1857
rect 2068 1857 2083 1895
rect 2090 1857 2105 1895
rect 2068 1855 2105 1857
rect 2107 1857 2116 1895
rect 2123 1857 2126 1895
rect 2107 1855 2126 1857
rect 1931 1811 1951 1813
rect 1931 1773 1934 1811
rect 1941 1773 1951 1811
rect 1953 1811 1990 1813
rect 1953 1773 1968 1811
rect 1975 1773 1990 1811
rect 1992 1811 2011 1813
rect 1992 1773 2001 1811
rect 2008 1773 2011 1811
rect 1475 1607 1525 1608
rect 1475 1604 1525 1605
rect 1482 1549 1522 1552
rect 1482 1542 1484 1549
rect 1482 1532 1522 1542
rect 1482 1515 1522 1530
rect 1482 1508 1484 1515
rect 1482 1493 1522 1508
rect 1482 1482 1522 1491
rect 1482 1475 1484 1482
rect 1482 1472 1522 1475
rect 1475 1434 1525 1435
rect 1741 1437 1791 1438
rect 1475 1431 1525 1432
rect 1741 1434 1791 1435
rect 1479 1372 1529 1373
rect 1744 1379 1784 1382
rect 1782 1372 1784 1379
rect 1479 1369 1529 1370
rect 1744 1362 1784 1372
rect 1744 1345 1784 1360
rect 1782 1338 1784 1345
rect 1744 1323 1784 1338
rect 1486 1314 1526 1317
rect 1486 1307 1488 1314
rect 1486 1297 1526 1307
rect 1486 1280 1526 1295
rect 1486 1273 1488 1280
rect 1486 1258 1526 1273
rect 1744 1312 1784 1321
rect 1782 1305 1784 1312
rect 1744 1302 1784 1305
rect 1741 1264 1791 1265
rect 1486 1247 1526 1256
rect 1486 1240 1488 1247
rect 1486 1237 1526 1240
rect 1741 1261 1791 1262
rect 1479 1199 1529 1200
rect 2230 1891 2233 1929
rect 2240 1891 2250 1929
rect 2252 1929 2289 1931
rect 2252 1891 2267 1929
rect 2274 1891 2289 1929
rect 2291 1929 2310 1931
rect 2291 1891 2300 1929
rect 2307 1891 2310 1929
rect 2230 1645 2233 1683
rect 2240 1645 2250 1683
rect 2230 1643 2250 1645
rect 2252 1645 2267 1683
rect 2274 1645 2289 1683
rect 2252 1643 2289 1645
rect 2291 1645 2300 1683
rect 2307 1645 2310 1683
rect 2291 1643 2310 1645
rect 2532 1646 2535 1684
rect 2542 1646 2552 1684
rect 2532 1644 2552 1646
rect 2554 1646 2569 1684
rect 2576 1646 2591 1684
rect 2554 1644 2591 1646
rect 2593 1646 2602 1684
rect 2609 1646 2612 1684
rect 2593 1644 2612 1646
rect 2230 1599 2250 1601
rect 2230 1561 2233 1599
rect 2240 1561 2250 1599
rect 2252 1599 2289 1601
rect 2252 1561 2267 1599
rect 2274 1561 2289 1599
rect 2291 1599 2310 1601
rect 2291 1561 2300 1599
rect 2307 1561 2310 1599
rect 2360 1559 2361 1609
rect 2363 1559 2364 1609
rect 2406 1600 2426 1602
rect 2406 1562 2409 1600
rect 2416 1562 2426 1600
rect 2428 1600 2465 1602
rect 2428 1562 2443 1600
rect 2450 1562 2465 1600
rect 2467 1600 2486 1602
rect 2467 1562 2476 1600
rect 2483 1562 2486 1600
rect 2532 1600 2552 1602
rect 2532 1562 2535 1600
rect 2542 1562 2552 1600
rect 2554 1600 2591 1602
rect 2554 1562 2569 1600
rect 2576 1562 2591 1600
rect 2593 1600 2612 1602
rect 2593 1562 2602 1600
rect 2609 1562 2612 1600
rect 2230 1315 2233 1353
rect 2240 1315 2250 1353
rect 2230 1313 2250 1315
rect 2252 1315 2267 1353
rect 2274 1315 2289 1353
rect 2252 1313 2289 1315
rect 2291 1315 2300 1353
rect 2307 1315 2310 1353
rect 2291 1313 2310 1315
rect 2230 1269 2250 1271
rect 2230 1231 2233 1269
rect 2240 1231 2250 1269
rect 2252 1269 2289 1271
rect 2252 1231 2267 1269
rect 2274 1231 2289 1269
rect 2291 1269 2310 1271
rect 2291 1231 2300 1269
rect 2307 1231 2310 1269
rect 1479 1196 1529 1197
rect 1732 1175 1782 1176
rect 1732 1172 1782 1173
rect 1735 1117 1775 1120
rect 1773 1110 1775 1117
rect 1735 1100 1775 1110
rect 1735 1083 1775 1098
rect 1773 1076 1775 1083
rect 1735 1061 1775 1076
rect 1735 1050 1775 1059
rect 1773 1043 1775 1050
rect 1735 1040 1775 1043
rect 1732 1002 1782 1003
rect 1732 999 1782 1000
rect 2230 985 2233 1023
rect 2240 985 2250 1023
rect 2230 983 2250 985
rect 2252 985 2267 1023
rect 2274 985 2289 1023
rect 2252 983 2289 985
rect 2291 985 2300 1023
rect 2307 985 2310 1023
rect 2291 983 2310 985
rect 2532 986 2535 1024
rect 2542 986 2552 1024
rect 2532 984 2552 986
rect 2554 986 2569 1024
rect 2576 986 2591 1024
rect 2554 984 2591 986
rect 2593 986 2602 1024
rect 2609 986 2612 1024
rect 2593 984 2612 986
rect 2230 939 2250 941
rect 2230 901 2233 939
rect 2240 901 2250 939
rect 2252 939 2289 941
rect 2252 901 2267 939
rect 2274 901 2289 939
rect 2291 939 2310 941
rect 2291 901 2300 939
rect 2307 901 2310 939
rect 2360 899 2361 949
rect 2363 899 2364 949
rect 2406 940 2426 942
rect 2406 902 2409 940
rect 2416 902 2426 940
rect 2428 940 2465 942
rect 2428 902 2443 940
rect 2450 902 2465 940
rect 2467 940 2486 942
rect 2467 902 2476 940
rect 2483 902 2486 940
rect 2532 940 2552 942
rect 2532 902 2535 940
rect 2542 902 2552 940
rect 2554 940 2591 942
rect 2554 902 2569 940
rect 2576 902 2591 940
rect 2593 940 2612 942
rect 2593 902 2602 940
rect 2609 902 2612 940
rect 2230 655 2233 693
rect 2240 655 2250 693
rect 2230 653 2250 655
rect 2252 655 2267 693
rect 2274 655 2289 693
rect 2252 653 2289 655
rect 2291 655 2300 693
rect 2307 655 2310 693
rect 2291 653 2310 655
rect 273 126 313 129
rect 311 119 313 126
rect 273 109 313 119
rect 355 126 395 129
rect 355 119 357 126
rect 273 92 313 107
rect 355 109 395 119
rect 311 85 313 92
rect 273 70 313 85
rect 355 92 395 107
rect 355 85 357 92
rect 355 70 395 85
rect 273 59 313 68
rect 311 52 313 59
rect 273 49 313 52
rect 355 59 395 68
rect 355 52 357 59
rect 355 49 395 52
<< ndcontact >>
rect 112 4252 150 4259
rect 186 4252 224 4259
rect 442 4252 480 4259
rect 516 4252 554 4259
rect 112 4186 150 4193
rect 186 4186 224 4193
rect 442 4186 480 4193
rect 516 4186 554 4193
rect 228 4132 248 4136
rect 228 4124 248 4128
rect 187 4076 225 4083
rect 187 4010 225 4017
rect 187 3950 225 3957
rect 443 3950 481 3957
rect 187 3884 225 3891
rect 443 3884 481 3891
rect 1140 3624 1160 3628
rect 1140 3616 1160 3620
rect 1099 3558 1137 3565
rect 1934 3546 1941 3584
rect 2000 3546 2007 3584
rect 112 3295 150 3302
rect 186 3295 224 3302
rect 442 3295 480 3302
rect 516 3295 554 3302
rect 1099 3492 1137 3499
rect 1140 3451 1160 3455
rect 1140 3443 1160 3447
rect 1099 3393 1137 3400
rect 1099 3327 1137 3334
rect 1141 3291 1161 3295
rect 1141 3283 1161 3287
rect 112 3229 150 3236
rect 186 3229 224 3236
rect 442 3229 480 3236
rect 516 3229 554 3236
rect 228 3175 248 3179
rect 228 3167 248 3171
rect 187 3119 225 3126
rect 187 3053 225 3060
rect 740 3188 747 3226
rect 806 3188 813 3226
rect 864 3189 871 3227
rect 930 3189 937 3227
rect 979 3189 986 3227
rect 1045 3189 1052 3227
rect 1810 3291 1817 3329
rect 1876 3291 1883 3329
rect 1934 3290 1941 3328
rect 2000 3290 2007 3328
rect 2233 3785 2240 3823
rect 2299 3785 2306 3823
rect 2233 3711 2240 3749
rect 2299 3711 2306 3749
rect 2535 3712 2542 3750
rect 2601 3712 2608 3750
rect 2356 3497 2360 3517
rect 2364 3497 2368 3517
rect 2233 3455 2240 3493
rect 2299 3455 2306 3493
rect 2409 3456 2416 3494
rect 2475 3456 2482 3494
rect 2233 3381 2240 3419
rect 2299 3381 2306 3419
rect 2535 3456 2542 3494
rect 2601 3456 2608 3494
rect 2049 3290 2056 3328
rect 2115 3290 2122 3328
rect 1108 3172 1146 3179
rect 187 2993 225 3000
rect 443 2993 481 3000
rect 187 2927 225 2934
rect 443 2927 481 2934
rect 112 2816 150 2823
rect 186 2816 224 2823
rect 442 2816 480 2823
rect 516 2816 554 2823
rect 112 2750 150 2757
rect 186 2750 224 2757
rect 442 2750 480 2757
rect 516 2750 554 2757
rect 228 2696 248 2700
rect 228 2688 248 2692
rect 187 2640 225 2647
rect 187 2574 225 2581
rect 864 2933 871 2971
rect 930 2933 937 2971
rect 811 2877 849 2884
rect 811 2811 849 2818
rect 787 2775 807 2779
rect 787 2767 807 2771
rect 1108 3106 1146 3113
rect 1150 3070 1170 3074
rect 1810 3068 1817 3106
rect 1876 3068 1883 3106
rect 1934 3069 1941 3107
rect 2000 3069 2007 3107
rect 2049 3069 2056 3107
rect 2115 3069 2122 3107
rect 1150 3062 1170 3066
rect 1109 2967 1147 2974
rect 1109 2901 1147 2908
rect 1151 2865 1171 2869
rect 1151 2857 1171 2861
rect 1151 2784 1171 2788
rect 1151 2776 1171 2780
rect 187 2514 225 2521
rect 443 2514 481 2521
rect 187 2448 225 2455
rect 443 2448 481 2455
rect 112 2337 150 2344
rect 186 2337 224 2344
rect 442 2337 480 2344
rect 516 2337 554 2344
rect 112 2271 150 2278
rect 186 2271 224 2278
rect 442 2271 480 2278
rect 516 2271 554 2278
rect 228 2217 248 2221
rect 228 2209 248 2213
rect 187 2161 225 2168
rect 187 2095 225 2102
rect 1110 2718 1148 2725
rect 1110 2652 1148 2659
rect 787 2646 807 2650
rect 787 2638 807 2642
rect 1151 2611 1171 2615
rect 811 2599 849 2606
rect 1151 2603 1171 2607
rect 811 2533 849 2540
rect 864 2446 871 2484
rect 930 2446 937 2484
rect 740 2191 747 2229
rect 806 2191 813 2229
rect 187 2035 225 2042
rect 443 2035 481 2042
rect 187 1969 225 1976
rect 443 1969 481 1976
rect 112 1858 150 1865
rect 186 1858 224 1865
rect 442 1858 480 1865
rect 516 1858 554 1865
rect 112 1792 150 1799
rect 186 1792 224 1799
rect 442 1792 480 1799
rect 516 1792 554 1799
rect 1199 2232 1203 2252
rect 1207 2232 1211 2252
rect 864 2190 871 2228
rect 930 2190 937 2228
rect 979 2190 986 2228
rect 1045 2190 1052 2228
rect 1094 2190 1101 2228
rect 1160 2190 1167 2228
rect 1934 2813 1941 2851
rect 2000 2813 2007 2851
rect 1387 2734 1407 2738
rect 1387 2726 1407 2730
rect 2233 3125 2240 3163
rect 2299 3125 2306 3163
rect 2233 3051 2240 3089
rect 2299 3051 2306 3089
rect 2535 3052 2542 3090
rect 2601 3052 2608 3090
rect 2356 2837 2360 2857
rect 2364 2837 2368 2857
rect 2233 2795 2240 2833
rect 2299 2795 2306 2833
rect 2409 2796 2416 2834
rect 2475 2796 2482 2834
rect 2233 2721 2240 2759
rect 2299 2721 2306 2759
rect 1410 2668 1448 2675
rect 2535 2796 2542 2834
rect 2601 2796 2608 2834
rect 1410 2602 1448 2609
rect 1387 2561 1407 2565
rect 1387 2553 1407 2557
rect 228 1738 248 1742
rect 228 1730 248 1734
rect 187 1682 225 1689
rect 187 1616 225 1623
rect 1094 2116 1101 2154
rect 1160 2116 1167 2154
rect 740 2062 747 2100
rect 806 2062 813 2100
rect 864 2063 871 2101
rect 930 2063 937 2101
rect 979 2063 986 2101
rect 1045 2063 1052 2101
rect 1199 2092 1203 2112
rect 1207 2092 1211 2112
rect 187 1556 225 1563
rect 443 1556 481 1563
rect 187 1490 225 1497
rect 443 1490 481 1497
rect 112 1379 150 1386
rect 186 1379 224 1386
rect 442 1379 480 1386
rect 516 1379 554 1386
rect 112 1313 150 1320
rect 186 1313 224 1320
rect 442 1313 480 1320
rect 516 1313 554 1320
rect 228 1259 248 1263
rect 228 1251 248 1255
rect 187 1203 225 1210
rect 187 1137 225 1144
rect 864 1807 871 1845
rect 930 1807 937 1845
rect 811 1751 849 1758
rect 811 1685 849 1692
rect 787 1649 807 1653
rect 787 1641 807 1645
rect 187 1077 225 1084
rect 443 1077 481 1084
rect 187 1011 225 1018
rect 443 1011 481 1018
rect 112 900 150 907
rect 186 900 224 907
rect 442 900 480 907
rect 516 900 554 907
rect 112 834 150 841
rect 186 834 224 841
rect 442 834 480 841
rect 516 834 554 841
rect 228 780 248 784
rect 228 772 248 776
rect 187 724 225 731
rect 187 658 225 665
rect 187 598 225 605
rect 443 598 481 605
rect 187 532 225 539
rect 443 532 481 539
rect 112 421 150 428
rect 186 421 224 428
rect 442 421 480 428
rect 516 421 554 428
rect 112 355 150 362
rect 186 355 224 362
rect 442 355 480 362
rect 516 355 554 362
rect 228 301 248 305
rect 228 293 248 297
rect 187 245 225 252
rect 187 179 225 186
rect 1934 2420 1941 2458
rect 2000 2420 2007 2458
rect 1450 2379 1470 2383
rect 1450 2371 1470 2375
rect 1473 2313 1511 2320
rect 1473 2247 1511 2254
rect 1450 2206 1470 2210
rect 1602 2209 1622 2213
rect 1450 2198 1470 2202
rect 1602 2201 1622 2205
rect 1454 2144 1474 2148
rect 1561 2143 1599 2150
rect 1454 2136 1474 2140
rect 1477 2078 1515 2085
rect 1561 2077 1599 2084
rect 1810 2165 1817 2203
rect 1876 2165 1883 2203
rect 1934 2164 1941 2202
rect 2000 2164 2007 2202
rect 2049 2164 2056 2202
rect 2115 2164 2122 2202
rect 1602 2036 1622 2040
rect 1602 2028 1622 2032
rect 1477 2012 1515 2019
rect 1199 1886 1203 1906
rect 1207 1886 1211 1906
rect 1094 1844 1101 1882
rect 1160 1844 1167 1882
rect 2233 2465 2240 2503
rect 2299 2465 2306 2503
rect 2233 2391 2240 2429
rect 2299 2391 2306 2429
rect 2535 2392 2542 2430
rect 2601 2392 2608 2430
rect 2356 2177 2360 2197
rect 2364 2177 2368 2197
rect 2233 2135 2240 2173
rect 2299 2135 2306 2173
rect 2409 2136 2416 2174
rect 2475 2136 2482 2174
rect 2233 2061 2240 2099
rect 2299 2061 2306 2099
rect 2535 2136 2542 2174
rect 2601 2136 2608 2174
rect 1454 1971 1474 1975
rect 1091 1733 1098 1771
rect 1157 1733 1164 1771
rect 1196 1709 1200 1729
rect 1204 1709 1208 1729
rect 1454 1963 1474 1967
rect 1810 1942 1817 1980
rect 1876 1942 1883 1980
rect 1934 1943 1941 1981
rect 2000 1943 2007 1981
rect 2049 1943 2056 1981
rect 2115 1943 2122 1981
rect 1087 1532 1094 1570
rect 1153 1532 1160 1570
rect 1192 1508 1196 1528
rect 1200 1508 1204 1528
rect 1192 1304 1196 1324
rect 1200 1304 1204 1324
rect 1087 1262 1094 1300
rect 1153 1262 1160 1300
rect 1087 1159 1094 1197
rect 1153 1159 1160 1197
rect 1192 1135 1196 1155
rect 1200 1135 1204 1155
rect 1934 1687 1941 1725
rect 2000 1687 2007 1725
rect 1547 1608 1567 1612
rect 1547 1600 1567 1604
rect 1570 1542 1608 1549
rect 1570 1476 1608 1483
rect 1547 1435 1567 1439
rect 1699 1438 1719 1442
rect 1547 1427 1567 1431
rect 1699 1430 1719 1434
rect 1551 1373 1571 1377
rect 1658 1372 1696 1379
rect 1551 1365 1571 1369
rect 1574 1307 1612 1314
rect 1658 1306 1696 1313
rect 1699 1265 1719 1269
rect 1699 1257 1719 1261
rect 1574 1241 1612 1248
rect 1551 1200 1571 1204
rect 2233 1805 2240 1843
rect 2299 1805 2306 1843
rect 2233 1731 2240 1769
rect 2299 1731 2306 1769
rect 2535 1732 2542 1770
rect 2601 1732 2608 1770
rect 2356 1517 2360 1537
rect 2364 1517 2368 1537
rect 2233 1475 2240 1513
rect 2299 1475 2306 1513
rect 2409 1476 2416 1514
rect 2475 1476 2482 1514
rect 2233 1401 2240 1439
rect 2299 1401 2306 1439
rect 2535 1476 2542 1514
rect 2601 1476 2608 1514
rect 1551 1192 1571 1196
rect 1690 1176 1710 1180
rect 1690 1168 1710 1172
rect 1649 1110 1687 1117
rect 1649 1044 1687 1051
rect 1690 1003 1710 1007
rect 1690 995 1710 999
rect 2233 1145 2240 1183
rect 2299 1145 2306 1183
rect 2233 1071 2240 1109
rect 2299 1071 2306 1109
rect 2535 1072 2542 1110
rect 2601 1072 2608 1110
rect 2356 857 2360 877
rect 2364 857 2368 877
rect 2233 815 2240 853
rect 2299 815 2306 853
rect 2409 816 2416 854
rect 2475 816 2482 854
rect 2233 741 2240 779
rect 2299 741 2306 779
rect 2535 816 2542 854
rect 2601 816 2608 854
rect 187 119 225 126
rect 443 119 481 126
rect 187 53 225 60
rect 443 53 481 60
<< pdcontact >>
rect 26 4252 64 4259
rect 272 4252 310 4259
rect 356 4252 394 4259
rect 26 4218 64 4225
rect 602 4252 640 4259
rect 272 4218 310 4225
rect 356 4218 394 4225
rect 602 4218 640 4225
rect 26 4185 64 4192
rect 272 4185 310 4192
rect 356 4185 394 4192
rect 602 4185 640 4192
rect 270 4132 320 4136
rect 270 4124 320 4128
rect 273 4076 311 4083
rect 273 4042 311 4049
rect 273 4009 311 4016
rect 273 3950 311 3957
rect 357 3950 395 3957
rect 273 3916 311 3923
rect 357 3916 395 3923
rect 273 3883 311 3890
rect 357 3883 395 3890
rect 2233 3871 2240 3909
rect 2267 3871 2274 3909
rect 2300 3871 2307 3909
rect 1182 3624 1232 3628
rect 1182 3616 1232 3620
rect 1185 3558 1223 3565
rect 1185 3524 1223 3531
rect 26 3295 64 3302
rect 272 3295 310 3302
rect 356 3295 394 3302
rect 26 3261 64 3268
rect 602 3295 640 3302
rect 272 3261 310 3268
rect 356 3261 394 3268
rect 1185 3491 1223 3498
rect 1182 3451 1232 3455
rect 1182 3443 1232 3447
rect 1934 3460 1941 3498
rect 1968 3460 1975 3498
rect 2001 3460 2008 3498
rect 1185 3393 1223 3400
rect 1185 3359 1223 3366
rect 1810 3377 1817 3415
rect 1844 3377 1851 3415
rect 1877 3377 1884 3415
rect 1185 3326 1223 3333
rect 1183 3291 1233 3295
rect 1183 3283 1233 3287
rect 602 3261 640 3268
rect 26 3228 64 3235
rect 272 3228 310 3235
rect 356 3228 394 3235
rect 602 3228 640 3235
rect 270 3175 320 3179
rect 270 3167 320 3171
rect 273 3119 311 3126
rect 273 3085 311 3092
rect 273 3052 311 3059
rect 1934 3376 1941 3414
rect 1968 3376 1975 3414
rect 2001 3376 2008 3414
rect 2049 3376 2056 3414
rect 2083 3376 2090 3414
rect 2116 3376 2123 3414
rect 2233 3625 2240 3663
rect 2267 3625 2274 3663
rect 2300 3625 2307 3663
rect 2535 3626 2542 3664
rect 2569 3626 2576 3664
rect 2602 3626 2609 3664
rect 2233 3541 2240 3579
rect 2267 3541 2274 3579
rect 2300 3541 2307 3579
rect 2356 3539 2360 3589
rect 2364 3539 2368 3589
rect 2409 3542 2416 3580
rect 2443 3542 2450 3580
rect 2476 3542 2483 3580
rect 2535 3542 2542 3580
rect 2569 3542 2576 3580
rect 2602 3542 2609 3580
rect 2233 3295 2240 3333
rect 2267 3295 2274 3333
rect 2300 3295 2307 3333
rect 2233 3211 2240 3249
rect 2267 3211 2274 3249
rect 2300 3211 2307 3249
rect 740 3102 747 3140
rect 774 3102 781 3140
rect 807 3102 814 3140
rect 1194 3172 1232 3179
rect 864 3103 871 3141
rect 898 3103 905 3141
rect 931 3103 938 3141
rect 979 3103 986 3141
rect 1013 3103 1020 3141
rect 1046 3103 1053 3141
rect 1194 3138 1232 3145
rect 864 3019 871 3057
rect 898 3019 905 3057
rect 931 3019 938 3057
rect 273 2993 311 3000
rect 357 2993 395 3000
rect 273 2959 311 2966
rect 357 2959 395 2966
rect 273 2926 311 2933
rect 357 2926 395 2933
rect 26 2816 64 2823
rect 272 2816 310 2823
rect 356 2816 394 2823
rect 26 2782 64 2789
rect 602 2816 640 2823
rect 272 2782 310 2789
rect 356 2782 394 2789
rect 602 2782 640 2789
rect 26 2749 64 2756
rect 272 2749 310 2756
rect 356 2749 394 2756
rect 602 2749 640 2756
rect 270 2696 320 2700
rect 270 2688 320 2692
rect 273 2640 311 2647
rect 273 2606 311 2613
rect 273 2573 311 2580
rect 725 2877 763 2884
rect 725 2843 763 2850
rect 725 2810 763 2817
rect 715 2775 765 2779
rect 715 2767 765 2771
rect 1194 3105 1232 3112
rect 1192 3070 1242 3074
rect 1192 3062 1242 3066
rect 1810 2982 1817 3020
rect 1844 2982 1851 3020
rect 1877 2982 1884 3020
rect 1195 2967 1233 2974
rect 1195 2933 1233 2940
rect 1195 2900 1233 2907
rect 1934 2983 1941 3021
rect 1968 2983 1975 3021
rect 2001 2983 2008 3021
rect 2049 2983 2056 3021
rect 2083 2983 2090 3021
rect 2116 2983 2123 3021
rect 1934 2899 1941 2937
rect 1968 2899 1975 2937
rect 2001 2899 2008 2937
rect 1193 2865 1243 2869
rect 1193 2857 1243 2861
rect 1193 2784 1243 2788
rect 1193 2776 1243 2780
rect 273 2514 311 2521
rect 357 2514 395 2521
rect 273 2480 311 2487
rect 357 2480 395 2487
rect 273 2447 311 2454
rect 357 2447 395 2454
rect 26 2337 64 2344
rect 272 2337 310 2344
rect 356 2337 394 2344
rect 26 2303 64 2310
rect 602 2337 640 2344
rect 272 2303 310 2310
rect 356 2303 394 2310
rect 602 2303 640 2310
rect 26 2270 64 2277
rect 272 2270 310 2277
rect 356 2270 394 2277
rect 602 2270 640 2277
rect 270 2217 320 2221
rect 270 2209 320 2213
rect 273 2161 311 2168
rect 273 2127 311 2134
rect 273 2094 311 2101
rect 1196 2718 1234 2725
rect 1196 2684 1234 2691
rect 715 2646 765 2650
rect 715 2638 765 2642
rect 1196 2651 1234 2658
rect 1193 2611 1243 2615
rect 725 2600 763 2607
rect 1193 2603 1243 2607
rect 725 2567 763 2574
rect 725 2533 763 2540
rect 740 2277 747 2315
rect 774 2277 781 2315
rect 807 2277 814 2315
rect 864 2360 871 2398
rect 898 2360 905 2398
rect 931 2360 938 2398
rect 864 2276 871 2314
rect 898 2276 905 2314
rect 931 2276 938 2314
rect 979 2276 986 2314
rect 1013 2276 1020 2314
rect 1046 2276 1053 2314
rect 1094 2276 1101 2314
rect 1128 2276 1135 2314
rect 1161 2276 1168 2314
rect 273 2035 311 2042
rect 357 2035 395 2042
rect 273 2001 311 2008
rect 357 2001 395 2008
rect 273 1968 311 1975
rect 357 1968 395 1975
rect 26 1858 64 1865
rect 272 1858 310 1865
rect 356 1858 394 1865
rect 26 1824 64 1831
rect 602 1858 640 1865
rect 272 1824 310 1831
rect 356 1824 394 1831
rect 602 1824 640 1831
rect 26 1791 64 1798
rect 272 1791 310 1798
rect 356 1791 394 1798
rect 1199 2274 1203 2324
rect 1207 2274 1211 2324
rect 1315 2734 1365 2738
rect 1315 2726 1365 2730
rect 2233 2965 2240 3003
rect 2267 2965 2274 3003
rect 2300 2965 2307 3003
rect 2535 2966 2542 3004
rect 2569 2966 2576 3004
rect 2602 2966 2609 3004
rect 2233 2881 2240 2919
rect 2267 2881 2274 2919
rect 2300 2881 2307 2919
rect 2356 2879 2360 2929
rect 2364 2879 2368 2929
rect 2409 2882 2416 2920
rect 2443 2882 2450 2920
rect 2476 2882 2483 2920
rect 2535 2882 2542 2920
rect 2569 2882 2576 2920
rect 2602 2882 2609 2920
rect 1324 2668 1362 2675
rect 1324 2634 1362 2641
rect 2233 2635 2240 2673
rect 2267 2635 2274 2673
rect 2300 2635 2307 2673
rect 1324 2601 1362 2608
rect 1315 2561 1365 2565
rect 1315 2553 1365 2557
rect 602 1791 640 1798
rect 270 1738 320 1742
rect 270 1730 320 1734
rect 273 1682 311 1689
rect 273 1648 311 1655
rect 273 1615 311 1622
rect 740 1976 747 2014
rect 774 1976 781 2014
rect 807 1976 814 2014
rect 864 1977 871 2015
rect 898 1977 905 2015
rect 931 1977 938 2015
rect 979 1977 986 2015
rect 1013 1977 1020 2015
rect 1046 1977 1053 2015
rect 864 1893 871 1931
rect 898 1893 905 1931
rect 931 1893 938 1931
rect 273 1556 311 1563
rect 357 1556 395 1563
rect 273 1522 311 1529
rect 357 1522 395 1529
rect 273 1489 311 1496
rect 357 1489 395 1496
rect 26 1379 64 1386
rect 272 1379 310 1386
rect 356 1379 394 1386
rect 26 1345 64 1352
rect 602 1379 640 1386
rect 272 1345 310 1352
rect 356 1345 394 1352
rect 602 1345 640 1352
rect 26 1312 64 1319
rect 272 1312 310 1319
rect 356 1312 394 1319
rect 602 1312 640 1319
rect 270 1259 320 1263
rect 270 1251 320 1255
rect 273 1203 311 1210
rect 273 1169 311 1176
rect 273 1136 311 1143
rect 725 1751 763 1758
rect 725 1717 763 1724
rect 725 1684 763 1691
rect 715 1649 765 1653
rect 715 1641 765 1645
rect 273 1077 311 1084
rect 357 1077 395 1084
rect 273 1043 311 1050
rect 357 1043 395 1050
rect 273 1010 311 1017
rect 357 1010 395 1017
rect 26 900 64 907
rect 272 900 310 907
rect 356 900 394 907
rect 26 866 64 873
rect 602 900 640 907
rect 272 866 310 873
rect 356 866 394 873
rect 602 866 640 873
rect 26 833 64 840
rect 272 833 310 840
rect 356 833 394 840
rect 602 833 640 840
rect 270 780 320 784
rect 270 772 320 776
rect 273 724 311 731
rect 273 690 311 697
rect 273 657 311 664
rect 273 598 311 605
rect 357 598 395 605
rect 273 564 311 571
rect 357 564 395 571
rect 273 531 311 538
rect 357 531 395 538
rect 26 421 64 428
rect 272 421 310 428
rect 356 421 394 428
rect 26 387 64 394
rect 602 421 640 428
rect 272 387 310 394
rect 356 387 394 394
rect 602 387 640 394
rect 26 354 64 361
rect 272 354 310 361
rect 356 354 394 361
rect 602 354 640 361
rect 270 301 320 305
rect 270 293 320 297
rect 273 245 311 252
rect 273 211 311 218
rect 273 178 311 185
rect 1094 2030 1101 2068
rect 1128 2030 1135 2068
rect 1161 2030 1168 2068
rect 1199 2020 1203 2070
rect 1207 2020 1211 2070
rect 2233 2551 2240 2589
rect 2267 2551 2274 2589
rect 2300 2551 2307 2589
rect 1378 2379 1428 2383
rect 1378 2371 1428 2375
rect 1387 2313 1425 2320
rect 1934 2334 1941 2372
rect 1968 2334 1975 2372
rect 2001 2334 2008 2372
rect 1387 2279 1425 2286
rect 1387 2246 1425 2253
rect 1810 2251 1817 2289
rect 1844 2251 1851 2289
rect 1877 2251 1884 2289
rect 1378 2206 1428 2210
rect 1644 2209 1694 2213
rect 1378 2198 1428 2202
rect 1644 2201 1694 2205
rect 1934 2250 1941 2288
rect 1968 2250 1975 2288
rect 2001 2250 2008 2288
rect 1382 2144 1432 2148
rect 1647 2143 1685 2150
rect 1382 2136 1432 2140
rect 1647 2109 1685 2116
rect 1391 2078 1429 2085
rect 1391 2044 1429 2051
rect 1647 2076 1685 2083
rect 2049 2250 2056 2288
rect 2083 2250 2090 2288
rect 2116 2250 2123 2288
rect 1644 2036 1694 2040
rect 1391 2011 1429 2018
rect 1644 2028 1694 2032
rect 1094 1930 1101 1968
rect 1128 1930 1135 1968
rect 1161 1930 1168 1968
rect 1199 1928 1203 1978
rect 1207 1928 1211 1978
rect 2233 2305 2240 2343
rect 2267 2305 2274 2343
rect 2300 2305 2307 2343
rect 2535 2306 2542 2344
rect 2569 2306 2576 2344
rect 2602 2306 2609 2344
rect 2233 2221 2240 2259
rect 2267 2221 2274 2259
rect 2300 2221 2307 2259
rect 2356 2219 2360 2269
rect 2364 2219 2368 2269
rect 2409 2222 2416 2260
rect 2443 2222 2450 2260
rect 2476 2222 2483 2260
rect 2535 2222 2542 2260
rect 2569 2222 2576 2260
rect 2602 2222 2609 2260
rect 1382 1971 1432 1975
rect 1382 1963 1432 1967
rect 1091 1647 1098 1685
rect 1125 1647 1132 1685
rect 1158 1647 1165 1685
rect 1196 1637 1200 1687
rect 1204 1637 1208 1687
rect 2233 1975 2240 2013
rect 2267 1975 2274 2013
rect 2300 1975 2307 2013
rect 1087 1446 1094 1484
rect 1121 1446 1128 1484
rect 1154 1446 1161 1484
rect 1192 1436 1196 1486
rect 1200 1436 1204 1486
rect 1087 1348 1094 1386
rect 1121 1348 1128 1386
rect 1154 1348 1161 1386
rect 1192 1346 1196 1396
rect 1200 1346 1204 1396
rect 1087 1073 1094 1111
rect 1121 1073 1128 1111
rect 1154 1073 1161 1111
rect 1192 1063 1196 1113
rect 1200 1063 1204 1113
rect 1810 1856 1817 1894
rect 1844 1856 1851 1894
rect 1877 1856 1884 1894
rect 1934 1857 1941 1895
rect 1968 1857 1975 1895
rect 2001 1857 2008 1895
rect 2049 1857 2056 1895
rect 2083 1857 2090 1895
rect 2116 1857 2123 1895
rect 1934 1773 1941 1811
rect 1968 1773 1975 1811
rect 2001 1773 2008 1811
rect 1475 1608 1525 1612
rect 1475 1600 1525 1604
rect 1484 1542 1522 1549
rect 1484 1508 1522 1515
rect 1484 1475 1522 1482
rect 1475 1435 1525 1439
rect 1741 1438 1791 1442
rect 1475 1427 1525 1431
rect 1741 1430 1791 1434
rect 1479 1373 1529 1377
rect 1744 1372 1782 1379
rect 1479 1365 1529 1369
rect 1744 1338 1782 1345
rect 1488 1307 1526 1314
rect 1488 1273 1526 1280
rect 1744 1305 1782 1312
rect 1741 1265 1791 1269
rect 1488 1240 1526 1247
rect 1741 1257 1791 1261
rect 1479 1200 1529 1204
rect 2233 1891 2240 1929
rect 2267 1891 2274 1929
rect 2300 1891 2307 1929
rect 2233 1645 2240 1683
rect 2267 1645 2274 1683
rect 2300 1645 2307 1683
rect 2535 1646 2542 1684
rect 2569 1646 2576 1684
rect 2602 1646 2609 1684
rect 2233 1561 2240 1599
rect 2267 1561 2274 1599
rect 2300 1561 2307 1599
rect 2356 1559 2360 1609
rect 2364 1559 2368 1609
rect 2409 1562 2416 1600
rect 2443 1562 2450 1600
rect 2476 1562 2483 1600
rect 2535 1562 2542 1600
rect 2569 1562 2576 1600
rect 2602 1562 2609 1600
rect 2233 1315 2240 1353
rect 2267 1315 2274 1353
rect 2300 1315 2307 1353
rect 2233 1231 2240 1269
rect 2267 1231 2274 1269
rect 2300 1231 2307 1269
rect 1479 1192 1529 1196
rect 1732 1176 1782 1180
rect 1732 1168 1782 1172
rect 1735 1110 1773 1117
rect 1735 1076 1773 1083
rect 1735 1043 1773 1050
rect 1732 1003 1782 1007
rect 1732 995 1782 999
rect 2233 985 2240 1023
rect 2267 985 2274 1023
rect 2300 985 2307 1023
rect 2535 986 2542 1024
rect 2569 986 2576 1024
rect 2602 986 2609 1024
rect 2233 901 2240 939
rect 2267 901 2274 939
rect 2300 901 2307 939
rect 2356 899 2360 949
rect 2364 899 2368 949
rect 2409 902 2416 940
rect 2443 902 2450 940
rect 2476 902 2483 940
rect 2535 902 2542 940
rect 2569 902 2576 940
rect 2602 902 2609 940
rect 2233 655 2240 693
rect 2267 655 2274 693
rect 2300 655 2307 693
rect 273 119 311 126
rect 357 119 395 126
rect 273 85 311 92
rect 357 85 395 92
rect 273 52 311 59
rect 357 52 395 59
<< psubstratepcontact >>
rect 165 4223 171 4231
rect 495 4223 501 4231
rect 166 4047 172 4055
rect 166 3921 172 3929
rect 496 3921 502 3929
rect 1078 3529 1084 3537
rect 1962 3599 1970 3605
rect 165 3266 171 3274
rect 495 3266 501 3274
rect 1078 3364 1084 3372
rect 166 3090 172 3098
rect 768 3241 776 3247
rect 892 3242 900 3248
rect 1007 3242 1015 3248
rect 1838 3270 1846 3276
rect 1962 3269 1970 3275
rect 2261 3764 2269 3770
rect 2563 3765 2571 3771
rect 2261 3434 2269 3440
rect 2437 3435 2445 3441
rect 2563 3435 2571 3441
rect 2077 3269 2085 3275
rect 1087 3143 1093 3151
rect 1838 3121 1846 3127
rect 166 2964 172 2972
rect 496 2964 502 2972
rect 165 2787 171 2795
rect 495 2787 501 2795
rect 166 2611 172 2619
rect 892 2912 900 2918
rect 864 2848 870 2856
rect 1962 3122 1970 3128
rect 2077 3122 2085 3128
rect 1088 2938 1094 2946
rect 166 2485 172 2493
rect 496 2485 502 2493
rect 165 2308 171 2316
rect 495 2308 501 2316
rect 166 2132 172 2140
rect 1089 2689 1095 2697
rect 864 2561 870 2569
rect 892 2499 900 2505
rect 768 2170 776 2176
rect 166 2006 172 2014
rect 496 2006 502 2014
rect 165 1829 171 1837
rect 495 1829 501 1837
rect 892 2169 900 2175
rect 1007 2169 1015 2175
rect 1122 2169 1130 2175
rect 1962 2792 1970 2798
rect 2261 3104 2269 3110
rect 2563 3105 2571 3111
rect 2261 2774 2269 2780
rect 2437 2775 2445 2781
rect 2563 2775 2571 2781
rect 1463 2639 1469 2647
rect 166 1653 172 1661
rect 768 2115 776 2121
rect 892 2116 900 2122
rect 1007 2116 1015 2122
rect 166 1527 172 1535
rect 496 1527 502 1535
rect 165 1350 171 1358
rect 495 1350 501 1358
rect 166 1174 172 1182
rect 892 1786 900 1792
rect 864 1722 870 1730
rect 166 1048 172 1056
rect 496 1048 502 1056
rect 165 871 171 879
rect 495 871 501 879
rect 166 695 172 703
rect 166 569 172 577
rect 496 569 502 577
rect 165 392 171 400
rect 495 392 501 400
rect 166 216 172 224
rect 1962 2473 1970 2479
rect 1526 2284 1532 2292
rect 1540 2114 1546 2122
rect 1838 2144 1846 2150
rect 1962 2143 1970 2149
rect 2077 2143 2085 2149
rect 1530 2049 1536 2057
rect 1838 1995 1846 2001
rect 1122 1823 1130 1829
rect 2261 2444 2269 2450
rect 2563 2445 2571 2451
rect 2261 2114 2269 2120
rect 2437 2115 2445 2121
rect 2563 2115 2571 2121
rect 1962 1996 1970 2002
rect 2077 1996 2085 2002
rect 1119 1786 1127 1792
rect 1115 1585 1123 1591
rect 1115 1241 1123 1247
rect 1115 1212 1123 1218
rect 1962 1666 1970 1672
rect 1623 1513 1629 1521
rect 1637 1343 1643 1351
rect 1627 1278 1633 1286
rect 2261 1784 2269 1790
rect 2563 1785 2571 1791
rect 2261 1454 2269 1460
rect 2437 1455 2445 1461
rect 2563 1455 2571 1461
rect 1628 1081 1634 1089
rect 2261 1124 2269 1130
rect 2563 1125 2571 1131
rect 2261 794 2269 800
rect 2437 795 2445 801
rect 2563 795 2571 801
rect 166 90 172 98
rect 496 90 502 98
<< nsubstratencontact >>
rect 0 4235 6 4243
rect 330 4235 336 4243
rect 660 4235 666 4243
rect 331 4059 337 4067
rect 331 3933 337 3941
rect 2249 3929 2257 3935
rect 1243 3541 1249 3549
rect 0 3278 6 3286
rect 330 3278 336 3286
rect 660 3278 666 3286
rect 1826 3435 1834 3441
rect 1243 3376 1249 3384
rect 331 3102 337 3110
rect 1950 3434 1958 3440
rect 2065 3434 2073 3440
rect 2249 3599 2257 3605
rect 2425 3600 2433 3606
rect 2551 3600 2559 3606
rect 2249 3269 2257 3275
rect 756 3076 764 3082
rect 1252 3155 1258 3163
rect 880 3077 888 3083
rect 331 2976 337 2984
rect 0 2799 6 2807
rect 330 2799 336 2807
rect 660 2799 666 2807
rect 331 2623 337 2631
rect 699 2860 705 2868
rect 995 3077 1003 3083
rect 1253 2950 1259 2958
rect 1826 2956 1834 2962
rect 1950 2957 1958 2963
rect 2065 2957 2073 2963
rect 331 2497 337 2505
rect 0 2320 6 2328
rect 330 2320 336 2328
rect 660 2320 666 2328
rect 331 2144 337 2152
rect 1254 2701 1260 2709
rect 699 2549 705 2557
rect 756 2335 764 2341
rect 880 2334 888 2340
rect 995 2334 1003 2340
rect 1110 2334 1118 2340
rect 331 2018 337 2026
rect 0 1841 6 1849
rect 330 1841 336 1849
rect 660 1841 666 1849
rect 2249 2939 2257 2945
rect 2425 2940 2433 2946
rect 2551 2940 2559 2946
rect 1298 2651 1304 2659
rect 2249 2609 2257 2615
rect 331 1665 337 1673
rect 756 1950 764 1956
rect 880 1951 888 1957
rect 331 1539 337 1547
rect 0 1362 6 1370
rect 330 1362 336 1370
rect 660 1362 666 1370
rect 331 1186 337 1194
rect 699 1734 705 1742
rect 331 1060 337 1068
rect 0 883 6 891
rect 330 883 336 891
rect 660 883 666 891
rect 331 707 337 715
rect 331 581 337 589
rect 0 404 6 412
rect 330 404 336 412
rect 660 404 666 412
rect 331 228 337 236
rect 995 1951 1003 1957
rect 1110 2004 1118 2010
rect 1110 1988 1118 1994
rect 1361 2296 1367 2304
rect 1826 2309 1834 2315
rect 1950 2308 1958 2314
rect 1705 2126 1711 2134
rect 1365 2061 1371 2069
rect 2065 2308 2073 2314
rect 2249 2279 2257 2285
rect 2425 2280 2433 2286
rect 2551 2280 2559 2286
rect 1107 1621 1115 1627
rect 2249 1949 2257 1955
rect 1103 1420 1111 1426
rect 1103 1406 1111 1412
rect 1103 1047 1111 1053
rect 1826 1830 1834 1836
rect 1950 1831 1958 1837
rect 2065 1831 2073 1837
rect 1458 1525 1464 1533
rect 1802 1355 1808 1363
rect 1462 1290 1468 1298
rect 2249 1619 2257 1625
rect 2425 1620 2433 1626
rect 2551 1620 2559 1626
rect 2249 1289 2257 1295
rect 1793 1093 1799 1101
rect 2249 959 2257 965
rect 2425 960 2433 966
rect 2551 960 2559 966
rect 2249 629 2257 635
rect 331 102 337 110
<< polysilicon >>
rect 83 4275 577 4277
rect 83 4267 85 4275
rect 95 4242 97 4246
rect 325 4245 342 4247
rect 325 4242 327 4245
rect 21 4240 24 4242
rect 64 4240 112 4242
rect 152 4240 155 4242
rect 181 4240 184 4242
rect 224 4240 272 4242
rect 312 4240 327 4242
rect 340 4242 342 4245
rect 575 4242 577 4275
rect 340 4240 354 4242
rect 394 4240 442 4242
rect 482 4240 485 4242
rect 511 4240 514 4242
rect 554 4240 602 4242
rect 642 4240 645 4242
rect 21 4201 24 4203
rect 64 4201 112 4203
rect 152 4201 155 4203
rect 181 4201 184 4203
rect 224 4201 272 4203
rect 312 4201 326 4203
rect 351 4201 354 4203
rect 394 4201 442 4203
rect 482 4201 490 4203
rect 511 4201 514 4203
rect 554 4201 602 4203
rect 642 4201 645 4203
rect 100 3984 102 4201
rect 324 4160 326 4201
rect 488 4172 490 4201
rect 488 4170 579 4172
rect 324 4158 348 4160
rect 590 4160 592 4201
rect 478 4158 592 4160
rect 225 4129 228 4131
rect 248 4129 270 4131
rect 320 4129 323 4131
rect 253 4066 255 4071
rect 182 4064 185 4066
rect 225 4064 273 4066
rect 313 4064 316 4066
rect 175 4025 185 4027
rect 225 4025 273 4027
rect 313 4025 316 4027
rect 175 4024 177 4025
rect 122 4022 177 4024
rect 436 3987 692 3989
rect 100 3982 188 3984
rect 252 3940 254 3944
rect 182 3938 185 3940
rect 225 3938 273 3940
rect 313 3938 316 3940
rect 412 3940 414 3946
rect 352 3938 355 3940
rect 395 3938 443 3940
rect 483 3938 486 3940
rect 182 3899 185 3901
rect 225 3899 273 3901
rect 313 3899 316 3901
rect 341 3899 355 3901
rect 395 3899 443 3901
rect 483 3899 486 3901
rect 237 3850 239 3899
rect 341 3861 343 3899
rect 308 3859 343 3861
rect 414 3850 416 3855
rect 237 3848 416 3850
rect 176 3762 181 3764
rect 690 3511 692 3987
rect 2250 3911 2252 3914
rect 2289 3911 2291 3914
rect 2250 3846 2252 3871
rect 2215 3844 2252 3846
rect 1137 3621 1140 3623
rect 1160 3621 1182 3623
rect 1232 3621 1235 3623
rect 1841 3610 2034 3612
rect 1181 3592 1301 3594
rect 1164 3548 1166 3554
rect 1094 3546 1097 3548
rect 1137 3546 1185 3548
rect 1225 3546 1228 3548
rect 436 3509 667 3511
rect 690 3509 777 3511
rect 1299 3545 1301 3592
rect 1841 3545 1843 3610
rect 1951 3586 1953 3589
rect 1990 3586 1992 3589
rect 1299 3543 1843 3545
rect 1951 3516 1953 3546
rect 1847 3514 1953 3516
rect 665 3493 667 3509
rect 1094 3507 1097 3509
rect 1137 3507 1185 3509
rect 1225 3507 1228 3509
rect 665 3491 688 3493
rect 83 3318 577 3320
rect 83 3310 85 3318
rect 95 3285 97 3289
rect 325 3288 342 3290
rect 325 3285 327 3288
rect 21 3283 24 3285
rect 64 3283 112 3285
rect 152 3283 155 3285
rect 181 3283 184 3285
rect 224 3283 272 3285
rect 312 3283 327 3285
rect 340 3285 342 3288
rect 575 3285 577 3318
rect 340 3283 354 3285
rect 394 3283 442 3285
rect 482 3283 485 3285
rect 511 3283 514 3285
rect 554 3283 602 3285
rect 642 3283 645 3285
rect 686 3273 688 3491
rect 1173 3476 1175 3507
rect 1168 3474 1175 3476
rect 1137 3448 1140 3450
rect 1160 3448 1182 3450
rect 1232 3448 1235 3450
rect 1164 3427 1166 3448
rect 1847 3431 1849 3514
rect 1951 3498 1953 3514
rect 1990 3498 1992 3546
rect 1951 3455 1953 3458
rect 1990 3447 1992 3458
rect 1827 3429 1849 3431
rect 1910 3445 1992 3447
rect 1164 3425 1264 3427
rect 1827 3417 1829 3429
rect 1866 3417 1868 3420
rect 1238 3387 1781 3389
rect 1238 3383 1240 3387
rect 1071 3381 1097 3383
rect 1137 3381 1185 3383
rect 1225 3381 1240 3383
rect 831 3273 833 3363
rect 1779 3356 1781 3387
rect 1827 3356 1829 3377
rect 1779 3354 1829 3356
rect 1090 3342 1097 3344
rect 1137 3342 1185 3344
rect 1225 3342 1725 3344
rect 1090 3282 1092 3342
rect 1138 3288 1141 3290
rect 1161 3288 1183 3290
rect 1233 3288 1236 3290
rect 686 3271 833 3273
rect 960 3280 1092 3282
rect 960 3260 962 3280
rect 686 3258 962 3260
rect 21 3244 24 3246
rect 64 3244 112 3246
rect 152 3244 155 3246
rect 181 3244 184 3246
rect 224 3244 272 3246
rect 312 3244 326 3246
rect 351 3244 354 3246
rect 394 3244 442 3246
rect 482 3244 490 3246
rect 511 3244 514 3246
rect 554 3244 602 3246
rect 642 3244 645 3246
rect 100 3027 102 3244
rect 324 3203 326 3244
rect 488 3215 490 3244
rect 488 3213 579 3215
rect 324 3201 348 3203
rect 590 3203 592 3244
rect 478 3201 592 3203
rect 225 3172 228 3174
rect 248 3172 270 3174
rect 320 3172 323 3174
rect 253 3109 255 3114
rect 182 3107 185 3109
rect 225 3107 273 3109
rect 313 3107 316 3109
rect 175 3068 185 3070
rect 225 3068 273 3070
rect 313 3068 316 3070
rect 175 3067 177 3068
rect 122 3065 177 3067
rect 686 3032 688 3258
rect 757 3228 759 3231
rect 796 3228 798 3231
rect 881 3229 883 3232
rect 920 3229 922 3232
rect 996 3229 998 3232
rect 1035 3229 1037 3232
rect 1723 3209 1725 3342
rect 1827 3329 1829 3354
rect 1866 3339 1868 3377
rect 1910 3361 1912 3445
rect 1951 3416 1953 3419
rect 1990 3416 1992 3419
rect 1951 3339 1953 3376
rect 1990 3348 1992 3376
rect 1984 3346 1992 3348
rect 1866 3337 1953 3339
rect 1866 3329 1868 3337
rect 1951 3328 1953 3337
rect 1990 3328 1992 3346
rect 1827 3285 1829 3289
rect 1866 3209 1868 3289
rect 1951 3285 1953 3288
rect 1990 3285 1992 3288
rect 1723 3207 1868 3209
rect 2032 3190 2034 3610
rect 2100 3516 2107 3518
rect 2066 3416 2068 3419
rect 2105 3416 2107 3516
rect 2066 3357 2068 3376
rect 2058 3355 2068 3357
rect 2066 3328 2068 3355
rect 2105 3328 2107 3376
rect 2140 3356 2172 3358
rect 2170 3345 2172 3356
rect 2215 3354 2217 3844
rect 2250 3823 2252 3844
rect 2289 3861 2291 3871
rect 2289 3859 2334 3861
rect 2289 3823 2291 3859
rect 2250 3780 2252 3783
rect 2289 3780 2291 3783
rect 2320 3759 2322 3848
rect 2289 3757 2322 3759
rect 2250 3751 2252 3754
rect 2289 3751 2291 3757
rect 2332 3747 2334 3859
rect 2552 3752 2554 3755
rect 2591 3752 2593 3755
rect 2250 3663 2252 3711
rect 2289 3663 2291 3711
rect 2552 3683 2554 3712
rect 2546 3681 2554 3683
rect 2552 3664 2554 3681
rect 2591 3664 2593 3712
rect 2637 3683 2644 3685
rect 2250 3611 2252 3623
rect 2289 3620 2291 3623
rect 2552 3621 2554 3624
rect 2245 3609 2252 3611
rect 2245 3596 2247 3609
rect 2245 3594 2252 3596
rect 2332 3595 2334 3617
rect 2591 3612 2593 3624
rect 2591 3610 2633 3612
rect 2250 3581 2252 3594
rect 2289 3593 2334 3595
rect 2289 3581 2291 3593
rect 2361 3589 2363 3592
rect 2250 3493 2252 3541
rect 2289 3493 2291 3541
rect 2426 3582 2428 3585
rect 2465 3582 2467 3585
rect 2552 3582 2554 3585
rect 2591 3582 2593 3585
rect 2631 3577 2633 3610
rect 2361 3517 2363 3539
rect 2426 3524 2428 3542
rect 2421 3522 2428 3524
rect 2361 3494 2363 3497
rect 2426 3494 2428 3522
rect 2465 3494 2467 3542
rect 2552 3523 2554 3542
rect 2548 3521 2554 3523
rect 2552 3494 2554 3521
rect 2591 3508 2593 3542
rect 2642 3508 2644 3683
rect 2591 3506 2644 3508
rect 2591 3494 2593 3506
rect 2250 3450 2252 3453
rect 2289 3450 2291 3453
rect 2426 3451 2428 3454
rect 2465 3446 2467 3454
rect 2465 3444 2470 3446
rect 2250 3421 2252 3424
rect 2289 3421 2291 3424
rect 2468 3391 2470 3444
rect 2215 3352 2225 3354
rect 2250 3345 2252 3381
rect 2170 3343 2252 3345
rect 2250 3333 2252 3343
rect 2289 3371 2291 3381
rect 2508 3371 2510 3457
rect 2552 3451 2554 3454
rect 2591 3451 2593 3454
rect 2289 3369 2510 3371
rect 2289 3333 2291 3369
rect 2250 3290 2252 3293
rect 2289 3290 2291 3293
rect 2066 3285 2068 3288
rect 2105 3285 2107 3288
rect 2250 3251 2252 3254
rect 2289 3251 2291 3254
rect 757 3140 759 3188
rect 796 3180 798 3188
rect 881 3180 883 3189
rect 796 3178 883 3180
rect 796 3140 798 3178
rect 757 3088 759 3100
rect 796 3097 798 3100
rect 757 3086 779 3088
rect 436 3030 688 3032
rect 100 3025 188 3027
rect 777 3003 779 3086
rect 831 3049 833 3178
rect 840 3072 842 3156
rect 881 3141 883 3178
rect 920 3171 922 3189
rect 914 3169 922 3171
rect 920 3141 922 3169
rect 996 3162 998 3189
rect 988 3160 998 3162
rect 996 3141 998 3160
rect 1035 3141 1037 3189
rect 1866 3188 2034 3190
rect 1071 3160 1081 3162
rect 1103 3160 1106 3162
rect 1146 3160 1194 3162
rect 1234 3160 1237 3162
rect 1079 3123 1081 3160
rect 1079 3121 1106 3123
rect 1146 3121 1194 3123
rect 1234 3121 1746 3123
rect 881 3089 883 3101
rect 920 3098 922 3101
rect 996 3098 998 3101
rect 881 3087 962 3089
rect 840 3070 922 3072
rect 881 3059 883 3062
rect 920 3059 922 3070
rect 881 3003 883 3019
rect 252 2983 254 2987
rect 777 3001 883 3003
rect 182 2981 185 2983
rect 225 2981 273 2983
rect 313 2981 316 2983
rect 412 2983 414 2989
rect 352 2981 355 2983
rect 395 2981 443 2983
rect 483 2981 486 2983
rect 792 2963 794 3001
rect 881 2971 883 3001
rect 920 2971 922 3019
rect 676 2961 794 2963
rect 182 2942 185 2944
rect 225 2942 273 2944
rect 313 2942 316 2944
rect 341 2942 355 2944
rect 395 2942 443 2944
rect 483 2942 486 2944
rect 237 2893 239 2942
rect 341 2904 343 2942
rect 308 2902 343 2904
rect 414 2893 416 2898
rect 237 2891 416 2893
rect 83 2839 577 2841
rect 83 2831 85 2839
rect 95 2806 97 2810
rect 325 2809 342 2811
rect 325 2806 327 2809
rect 21 2804 24 2806
rect 64 2804 112 2806
rect 152 2804 155 2806
rect 181 2804 184 2806
rect 224 2804 272 2806
rect 312 2804 327 2806
rect 340 2806 342 2809
rect 575 2806 577 2839
rect 340 2804 354 2806
rect 394 2804 442 2806
rect 482 2804 485 2806
rect 511 2804 514 2806
rect 554 2804 602 2806
rect 642 2804 645 2806
rect 21 2765 24 2767
rect 64 2765 112 2767
rect 152 2765 155 2767
rect 181 2765 184 2767
rect 224 2765 272 2767
rect 312 2765 326 2767
rect 351 2765 354 2767
rect 394 2765 442 2767
rect 482 2765 490 2767
rect 511 2765 514 2767
rect 554 2765 602 2767
rect 642 2765 645 2767
rect 100 2548 102 2765
rect 324 2724 326 2765
rect 488 2736 490 2765
rect 488 2734 579 2736
rect 324 2722 348 2724
rect 590 2724 592 2765
rect 478 2722 592 2724
rect 225 2693 228 2695
rect 248 2693 270 2695
rect 320 2693 323 2695
rect 253 2630 255 2635
rect 182 2628 185 2630
rect 225 2628 273 2630
rect 313 2628 316 2630
rect 175 2589 185 2591
rect 225 2589 273 2591
rect 313 2589 316 2591
rect 175 2588 177 2589
rect 122 2586 177 2588
rect 676 2553 678 2961
rect 792 2867 794 2961
rect 881 2928 883 2931
rect 920 2928 922 2931
rect 720 2865 723 2867
rect 763 2865 811 2867
rect 851 2865 854 2867
rect 794 2828 796 2832
rect 720 2826 723 2828
rect 763 2826 811 2828
rect 851 2826 854 2828
rect 712 2772 715 2774
rect 765 2772 787 2774
rect 807 2772 810 2774
rect 960 2746 962 3087
rect 1035 3001 1037 3101
rect 1030 2999 1037 3001
rect 1079 2918 1081 3121
rect 1744 3114 1746 3121
rect 1744 3112 1829 3114
rect 1827 3108 1829 3112
rect 1866 3108 1868 3188
rect 2250 3186 2252 3211
rect 2215 3184 2252 3186
rect 1951 3109 1953 3112
rect 1990 3109 1992 3112
rect 2066 3109 2068 3112
rect 2105 3109 2107 3112
rect 1147 3067 1150 3069
rect 1170 3067 1192 3069
rect 1242 3067 1245 3069
rect 1827 3020 1829 3068
rect 1866 3060 1868 3068
rect 1951 3060 1953 3069
rect 1866 3058 1953 3060
rect 1866 3020 1868 3058
rect 1168 3001 1285 3003
rect 1168 2957 1170 3001
rect 1827 2968 1829 2980
rect 1866 2977 1868 2980
rect 1827 2966 1849 2968
rect 1088 2955 1107 2957
rect 1147 2955 1195 2957
rect 1235 2955 1238 2957
rect 1079 2916 1107 2918
rect 1147 2916 1195 2918
rect 1235 2916 1238 2918
rect 1847 2883 1849 2966
rect 1910 2952 1912 3036
rect 1951 3021 1953 3058
rect 1990 3051 1992 3069
rect 1984 3049 1992 3051
rect 1990 3021 1992 3049
rect 2066 3042 2068 3069
rect 2058 3040 2068 3042
rect 2066 3021 2068 3040
rect 2105 3021 2107 3069
rect 2144 3040 2172 3042
rect 1951 2978 1953 2981
rect 1990 2978 1992 2981
rect 2066 2978 2068 2981
rect 1910 2950 1992 2952
rect 1951 2939 1953 2942
rect 1990 2939 1992 2950
rect 1951 2883 1953 2899
rect 1847 2881 1953 2883
rect 1148 2862 1151 2864
rect 1171 2862 1193 2864
rect 1243 2862 1246 2864
rect 1951 2851 1953 2881
rect 1990 2851 1992 2899
rect 2105 2881 2107 2981
rect 2100 2879 2107 2881
rect 1229 2827 1274 2829
rect 1148 2781 1151 2783
rect 1171 2781 1193 2783
rect 1243 2781 1246 2783
rect 436 2551 678 2553
rect 691 2744 962 2746
rect 100 2546 188 2548
rect 252 2504 254 2508
rect 182 2502 185 2504
rect 225 2502 273 2504
rect 313 2502 316 2504
rect 412 2504 414 2510
rect 352 2502 355 2504
rect 395 2502 443 2504
rect 483 2502 486 2504
rect 182 2463 185 2465
rect 225 2463 273 2465
rect 313 2463 316 2465
rect 341 2463 355 2465
rect 395 2463 443 2465
rect 483 2463 486 2465
rect 237 2414 239 2463
rect 341 2425 343 2463
rect 308 2423 343 2425
rect 414 2414 416 2419
rect 237 2412 416 2414
rect 83 2360 577 2362
rect 83 2352 85 2360
rect 95 2327 97 2331
rect 325 2330 342 2332
rect 325 2327 327 2330
rect 21 2325 24 2327
rect 64 2325 112 2327
rect 152 2325 155 2327
rect 181 2325 184 2327
rect 224 2325 272 2327
rect 312 2325 327 2327
rect 340 2327 342 2330
rect 575 2327 577 2360
rect 340 2325 354 2327
rect 394 2325 442 2327
rect 482 2325 485 2327
rect 511 2325 514 2327
rect 554 2325 602 2327
rect 642 2325 645 2327
rect 21 2286 24 2288
rect 64 2286 112 2288
rect 152 2286 155 2288
rect 181 2286 184 2288
rect 224 2286 272 2288
rect 312 2286 326 2288
rect 351 2286 354 2288
rect 394 2286 442 2288
rect 482 2286 490 2288
rect 511 2286 514 2288
rect 554 2286 602 2288
rect 642 2286 645 2288
rect 100 2069 102 2286
rect 324 2245 326 2286
rect 488 2257 490 2286
rect 488 2255 579 2257
rect 324 2243 348 2245
rect 590 2245 592 2286
rect 478 2243 592 2245
rect 225 2214 228 2216
rect 248 2214 270 2216
rect 320 2214 323 2216
rect 253 2151 255 2156
rect 182 2149 185 2151
rect 225 2149 273 2151
rect 313 2149 316 2151
rect 175 2110 185 2112
rect 225 2110 273 2112
rect 313 2110 316 2112
rect 175 2109 177 2110
rect 122 2107 177 2109
rect 691 2074 693 2744
rect 1175 2708 1177 2714
rect 1105 2706 1108 2708
rect 1148 2706 1196 2708
rect 1236 2706 1239 2708
rect 1105 2667 1108 2669
rect 1148 2667 1196 2669
rect 1236 2667 1239 2669
rect 712 2643 715 2645
rect 765 2643 787 2645
rect 807 2643 810 2645
rect 1184 2636 1186 2667
rect 1179 2634 1186 2636
rect 1148 2608 1151 2610
rect 1171 2608 1193 2610
rect 1243 2608 1246 2610
rect 720 2589 723 2591
rect 763 2589 811 2591
rect 851 2589 854 2591
rect 794 2585 796 2589
rect 720 2550 723 2552
rect 763 2550 811 2552
rect 851 2550 854 2552
rect 792 2416 794 2550
rect 881 2486 883 2489
rect 920 2486 922 2489
rect 881 2416 883 2446
rect 777 2414 883 2416
rect 777 2331 779 2414
rect 881 2398 883 2414
rect 920 2398 922 2446
rect 1030 2416 1037 2418
rect 757 2329 779 2331
rect 757 2317 759 2329
rect 796 2317 798 2320
rect 757 2229 759 2277
rect 796 2239 798 2277
rect 831 2239 833 2368
rect 881 2355 883 2358
rect 920 2347 922 2358
rect 840 2345 922 2347
rect 840 2261 842 2345
rect 881 2316 883 2319
rect 920 2316 922 2319
rect 996 2316 998 2319
rect 1035 2316 1037 2416
rect 1111 2316 1113 2319
rect 1150 2316 1152 2567
rect 1204 2324 1206 2327
rect 881 2239 883 2276
rect 920 2248 922 2276
rect 996 2257 998 2276
rect 988 2255 998 2257
rect 914 2246 922 2248
rect 796 2237 883 2239
rect 796 2229 798 2237
rect 757 2148 759 2189
rect 796 2186 798 2189
rect 436 2072 693 2074
rect 711 2146 759 2148
rect 100 2067 188 2069
rect 252 2025 254 2029
rect 182 2023 185 2025
rect 225 2023 273 2025
rect 313 2023 316 2025
rect 412 2025 414 2031
rect 352 2023 355 2025
rect 395 2023 443 2025
rect 483 2023 486 2025
rect 182 1984 185 1986
rect 225 1984 273 1986
rect 313 1984 316 1986
rect 341 1984 355 1986
rect 395 1984 443 1986
rect 483 1984 486 1986
rect 237 1935 239 1984
rect 341 1946 343 1984
rect 308 1944 343 1946
rect 414 1935 416 1940
rect 237 1933 416 1935
rect 83 1881 577 1883
rect 83 1873 85 1881
rect 95 1848 97 1852
rect 325 1851 342 1853
rect 325 1848 327 1851
rect 21 1846 24 1848
rect 64 1846 112 1848
rect 152 1846 155 1848
rect 181 1846 184 1848
rect 224 1846 272 1848
rect 312 1846 327 1848
rect 340 1848 342 1851
rect 575 1848 577 1881
rect 340 1846 354 1848
rect 394 1846 442 1848
rect 482 1846 485 1848
rect 511 1846 514 1848
rect 554 1846 602 1848
rect 642 1846 645 1848
rect 21 1807 24 1809
rect 64 1807 112 1809
rect 152 1807 155 1809
rect 181 1807 184 1809
rect 224 1807 272 1809
rect 312 1807 326 1809
rect 351 1807 354 1809
rect 394 1807 442 1809
rect 482 1807 490 1809
rect 511 1807 514 1809
rect 554 1807 602 1809
rect 642 1807 645 1809
rect 100 1590 102 1807
rect 324 1766 326 1807
rect 488 1778 490 1807
rect 488 1776 579 1778
rect 324 1764 348 1766
rect 590 1766 592 1807
rect 711 1806 713 2146
rect 831 2136 833 2237
rect 881 2228 883 2237
rect 920 2228 922 2246
rect 996 2228 998 2255
rect 1035 2228 1037 2276
rect 1111 2257 1113 2276
rect 1071 2255 1113 2257
rect 1111 2228 1113 2255
rect 1150 2228 1152 2276
rect 1204 2252 1206 2274
rect 1204 2229 1206 2232
rect 881 2185 883 2188
rect 920 2185 922 2188
rect 996 2185 998 2188
rect 1035 2185 1037 2188
rect 1111 2156 1113 2188
rect 1150 2185 1152 2188
rect 1272 2164 1274 2827
rect 1951 2808 1953 2811
rect 1990 2808 1992 2811
rect 1312 2731 1315 2733
rect 1365 2731 1387 2733
rect 1407 2731 1410 2733
rect 2170 2685 2172 3040
rect 2215 2694 2217 3184
rect 2250 3163 2252 3184
rect 2289 3201 2291 3211
rect 2289 3199 2334 3201
rect 2289 3163 2291 3199
rect 2250 3120 2252 3123
rect 2289 3120 2291 3123
rect 2320 3099 2322 3188
rect 2289 3097 2322 3099
rect 2250 3091 2252 3094
rect 2289 3091 2291 3097
rect 2332 3087 2334 3199
rect 2552 3092 2554 3095
rect 2591 3092 2593 3095
rect 2250 3003 2252 3051
rect 2289 3003 2291 3051
rect 2552 3023 2554 3052
rect 2546 3021 2554 3023
rect 2552 3004 2554 3021
rect 2591 3004 2593 3052
rect 2637 3023 2644 3025
rect 2250 2951 2252 2963
rect 2289 2960 2291 2963
rect 2552 2961 2554 2964
rect 2245 2949 2252 2951
rect 2245 2936 2247 2949
rect 2245 2934 2252 2936
rect 2332 2935 2334 2957
rect 2591 2952 2593 2964
rect 2591 2950 2633 2952
rect 2250 2921 2252 2934
rect 2289 2933 2334 2935
rect 2289 2921 2291 2933
rect 2361 2929 2363 2932
rect 2250 2833 2252 2881
rect 2289 2833 2291 2881
rect 2426 2922 2428 2925
rect 2465 2922 2467 2925
rect 2552 2922 2554 2925
rect 2591 2922 2593 2925
rect 2631 2917 2633 2950
rect 2361 2857 2363 2879
rect 2426 2864 2428 2882
rect 2421 2862 2428 2864
rect 2361 2834 2363 2837
rect 2426 2834 2428 2862
rect 2465 2834 2467 2882
rect 2552 2863 2554 2882
rect 2548 2861 2554 2863
rect 2552 2834 2554 2861
rect 2591 2848 2593 2882
rect 2642 2848 2644 3023
rect 2591 2846 2644 2848
rect 2591 2834 2593 2846
rect 2250 2790 2252 2793
rect 2289 2790 2291 2793
rect 2426 2791 2428 2794
rect 2465 2786 2467 2794
rect 2465 2784 2470 2786
rect 2250 2761 2252 2764
rect 2289 2761 2291 2764
rect 2468 2731 2470 2784
rect 2215 2692 2225 2694
rect 2250 2685 2252 2721
rect 2170 2683 2252 2685
rect 2250 2673 2252 2683
rect 2289 2711 2291 2721
rect 2508 2711 2510 2797
rect 2552 2791 2554 2794
rect 2591 2791 2593 2794
rect 2289 2709 2510 2711
rect 2289 2673 2291 2709
rect 1381 2658 1383 2664
rect 1319 2656 1322 2658
rect 1362 2656 1410 2658
rect 1450 2656 1453 2658
rect 2250 2630 2252 2633
rect 2289 2630 2291 2633
rect 1319 2617 1322 2619
rect 1362 2617 1410 2619
rect 1450 2617 1453 2619
rect 1372 2586 1374 2617
rect 1385 2594 1396 2596
rect 1394 2590 1396 2594
rect 2250 2591 2252 2594
rect 2289 2591 2291 2594
rect 1394 2588 1804 2590
rect 1372 2584 1379 2586
rect 1312 2558 1315 2560
rect 1365 2558 1387 2560
rect 1407 2558 1410 2560
rect 1150 2162 1274 2164
rect 1150 2156 1152 2162
rect 684 1804 713 1806
rect 719 2134 833 2136
rect 478 1764 592 1766
rect 225 1735 228 1737
rect 248 1735 270 1737
rect 320 1735 323 1737
rect 253 1672 255 1677
rect 182 1670 185 1672
rect 225 1670 273 1672
rect 313 1670 316 1672
rect 175 1631 185 1633
rect 225 1631 273 1633
rect 313 1631 316 1633
rect 175 1630 177 1631
rect 122 1628 177 1630
rect 684 1595 686 1804
rect 719 1788 721 2134
rect 757 2102 759 2105
rect 796 2102 798 2105
rect 881 2103 883 2106
rect 920 2103 922 2106
rect 996 2103 998 2106
rect 1035 2103 1037 2106
rect 1111 2068 1113 2116
rect 1150 2068 1152 2116
rect 1204 2112 1206 2115
rect 1204 2070 1206 2092
rect 757 2014 759 2062
rect 796 2054 798 2062
rect 881 2054 883 2063
rect 796 2052 883 2054
rect 796 2014 798 2052
rect 757 1962 759 1974
rect 796 1971 798 1974
rect 757 1960 779 1962
rect 777 1877 779 1960
rect 831 1923 833 2052
rect 840 1946 842 2030
rect 881 2015 883 2052
rect 920 2045 922 2063
rect 914 2043 922 2045
rect 920 2015 922 2043
rect 996 2036 998 2063
rect 988 2034 998 2036
rect 996 2015 998 2034
rect 1035 2015 1037 2063
rect 1071 2034 1077 2036
rect 881 1963 883 1975
rect 920 1972 922 1975
rect 996 1972 998 1975
rect 881 1961 959 1963
rect 840 1944 922 1946
rect 881 1933 883 1936
rect 920 1933 922 1944
rect 881 1877 883 1893
rect 777 1875 883 1877
rect 436 1593 686 1595
rect 692 1786 721 1788
rect 100 1588 188 1590
rect 252 1546 254 1550
rect 182 1544 185 1546
rect 225 1544 273 1546
rect 313 1544 316 1546
rect 412 1546 414 1552
rect 352 1544 355 1546
rect 395 1544 443 1546
rect 483 1544 486 1546
rect 182 1505 185 1507
rect 225 1505 273 1507
rect 313 1505 316 1507
rect 341 1505 355 1507
rect 395 1505 443 1507
rect 483 1505 486 1507
rect 237 1456 239 1505
rect 341 1467 343 1505
rect 308 1465 343 1467
rect 414 1456 416 1461
rect 237 1454 416 1456
rect 83 1402 577 1404
rect 83 1394 85 1402
rect 95 1369 97 1373
rect 325 1372 342 1374
rect 325 1369 327 1372
rect 21 1367 24 1369
rect 64 1367 112 1369
rect 152 1367 155 1369
rect 181 1367 184 1369
rect 224 1367 272 1369
rect 312 1367 327 1369
rect 340 1369 342 1372
rect 575 1369 577 1402
rect 340 1367 354 1369
rect 394 1367 442 1369
rect 482 1367 485 1369
rect 511 1367 514 1369
rect 554 1367 602 1369
rect 642 1367 645 1369
rect 21 1328 24 1330
rect 64 1328 112 1330
rect 152 1328 155 1330
rect 181 1328 184 1330
rect 224 1328 272 1330
rect 312 1328 326 1330
rect 351 1328 354 1330
rect 394 1328 442 1330
rect 482 1328 490 1330
rect 511 1328 514 1330
rect 554 1328 602 1330
rect 642 1328 645 1330
rect 100 1111 102 1328
rect 324 1287 326 1328
rect 488 1299 490 1328
rect 488 1297 579 1299
rect 324 1285 348 1287
rect 590 1287 592 1328
rect 478 1285 592 1287
rect 225 1256 228 1258
rect 248 1256 270 1258
rect 320 1256 323 1258
rect 253 1193 255 1198
rect 182 1191 185 1193
rect 225 1191 273 1193
rect 313 1191 316 1193
rect 175 1152 185 1154
rect 225 1152 273 1154
rect 313 1152 316 1154
rect 175 1151 177 1152
rect 122 1149 177 1151
rect 692 1116 694 1786
rect 792 1741 794 1875
rect 881 1845 883 1875
rect 920 1845 922 1893
rect 881 1802 883 1805
rect 920 1802 922 1805
rect 720 1739 723 1741
rect 763 1739 811 1741
rect 851 1739 882 1741
rect 794 1702 796 1706
rect 720 1700 723 1702
rect 763 1700 811 1702
rect 851 1700 854 1702
rect 712 1646 715 1648
rect 765 1646 787 1648
rect 807 1646 810 1648
rect 436 1114 694 1116
rect 100 1109 188 1111
rect 252 1067 254 1071
rect 182 1065 185 1067
rect 225 1065 273 1067
rect 313 1065 316 1067
rect 412 1067 414 1073
rect 352 1065 355 1067
rect 395 1065 443 1067
rect 483 1065 486 1067
rect 182 1026 185 1028
rect 225 1026 273 1028
rect 313 1026 316 1028
rect 341 1026 355 1028
rect 395 1026 443 1028
rect 483 1026 486 1028
rect 237 977 239 1026
rect 341 988 343 1026
rect 308 986 343 988
rect 414 977 416 982
rect 237 975 416 977
rect 83 923 577 925
rect 83 915 85 923
rect 95 890 97 894
rect 325 893 342 895
rect 325 890 327 893
rect 21 888 24 890
rect 64 888 112 890
rect 152 888 155 890
rect 181 888 184 890
rect 224 888 272 890
rect 312 888 327 890
rect 340 890 342 893
rect 575 890 577 923
rect 340 888 354 890
rect 394 888 442 890
rect 482 888 485 890
rect 511 888 514 890
rect 554 888 602 890
rect 642 888 645 890
rect 21 849 24 851
rect 64 849 112 851
rect 152 849 155 851
rect 181 849 184 851
rect 224 849 272 851
rect 312 849 326 851
rect 351 849 354 851
rect 394 849 442 851
rect 482 849 490 851
rect 511 849 514 851
rect 554 849 602 851
rect 642 849 645 851
rect 100 632 102 849
rect 324 808 326 849
rect 488 820 490 849
rect 488 818 579 820
rect 324 806 348 808
rect 590 808 592 849
rect 478 806 592 808
rect 225 777 228 779
rect 248 777 270 779
rect 320 777 323 779
rect 253 714 255 719
rect 182 712 185 714
rect 225 712 273 714
rect 313 712 316 714
rect 175 673 185 675
rect 225 673 273 675
rect 313 673 316 675
rect 175 672 177 673
rect 122 670 177 672
rect 880 637 882 1739
rect 436 635 882 637
rect 100 630 188 632
rect 252 588 254 592
rect 182 586 185 588
rect 225 586 273 588
rect 313 586 316 588
rect 412 588 414 594
rect 352 586 355 588
rect 395 586 443 588
rect 483 586 486 588
rect 182 547 185 549
rect 225 547 273 549
rect 313 547 316 549
rect 341 547 355 549
rect 395 547 443 549
rect 483 547 486 549
rect 237 498 239 547
rect 341 509 343 547
rect 308 507 343 509
rect 414 498 416 503
rect 237 496 416 498
rect 83 444 577 446
rect 83 436 85 444
rect 95 411 97 415
rect 325 414 342 416
rect 325 411 327 414
rect 21 409 24 411
rect 64 409 112 411
rect 152 409 155 411
rect 181 409 184 411
rect 224 409 272 411
rect 312 409 327 411
rect 340 411 342 414
rect 575 411 577 444
rect 340 409 354 411
rect 394 409 442 411
rect 482 409 485 411
rect 511 409 514 411
rect 554 409 602 411
rect 642 409 645 411
rect 21 370 24 372
rect 64 370 112 372
rect 152 370 155 372
rect 181 370 184 372
rect 224 370 272 372
rect 312 370 326 372
rect 351 370 354 372
rect 394 370 442 372
rect 482 370 490 372
rect 511 370 514 372
rect 554 370 602 372
rect 642 370 645 372
rect 100 153 102 370
rect 324 329 326 370
rect 488 341 490 370
rect 488 339 579 341
rect 324 327 348 329
rect 590 329 592 370
rect 478 327 592 329
rect 225 298 228 300
rect 248 298 270 300
rect 320 298 323 300
rect 253 235 255 240
rect 182 233 185 235
rect 225 233 273 235
rect 313 233 316 235
rect 175 194 185 196
rect 225 194 273 196
rect 313 194 316 196
rect 175 193 177 194
rect 122 191 177 193
rect 957 158 959 1961
rect 1035 1875 1037 1975
rect 1030 1873 1037 1875
rect 1075 1716 1077 2034
rect 1111 2016 1113 2028
rect 1150 2025 1152 2028
rect 1204 2017 1206 2020
rect 1111 2014 1126 2016
rect 1124 1984 1126 2014
rect 1307 2001 1309 2522
rect 1802 2507 1804 2588
rect 2250 2526 2252 2551
rect 2215 2524 2252 2526
rect 1802 2505 2028 2507
rect 1951 2460 1953 2463
rect 1990 2460 1992 2463
rect 1322 2406 1446 2408
rect 1444 2378 1446 2406
rect 1951 2390 1953 2420
rect 1847 2388 1953 2390
rect 1375 2376 1378 2378
rect 1428 2376 1450 2378
rect 1470 2376 1473 2378
rect 1444 2303 1446 2309
rect 1847 2305 1849 2388
rect 1951 2372 1953 2388
rect 1990 2372 1992 2420
rect 1951 2329 1953 2332
rect 1990 2321 1992 2332
rect 1827 2303 1849 2305
rect 1910 2319 1992 2321
rect 1382 2301 1385 2303
rect 1425 2301 1473 2303
rect 1513 2301 1516 2303
rect 1827 2291 1829 2303
rect 1866 2291 1868 2294
rect 1382 2262 1385 2264
rect 1425 2262 1473 2264
rect 1513 2262 1516 2264
rect 1435 2231 1437 2262
rect 1448 2239 1458 2241
rect 1435 2229 1442 2231
rect 1456 2229 1458 2239
rect 1545 2237 1628 2239
rect 1545 2229 1547 2237
rect 1456 2227 1547 2229
rect 1626 2208 1628 2237
rect 1599 2206 1602 2208
rect 1622 2206 1644 2208
rect 1694 2206 1697 2208
rect 1375 2203 1378 2205
rect 1428 2203 1450 2205
rect 1470 2203 1473 2205
rect 1444 2189 1446 2203
rect 1827 2203 1829 2251
rect 1866 2213 1868 2251
rect 1910 2235 1912 2319
rect 1951 2290 1953 2293
rect 1990 2290 1992 2293
rect 1951 2213 1953 2250
rect 1990 2222 1992 2250
rect 1984 2220 1992 2222
rect 1866 2211 1953 2213
rect 1866 2203 1868 2211
rect 1314 2187 1446 2189
rect 1314 2179 1316 2187
rect 1345 2180 1535 2182
rect 1111 1982 1126 1984
rect 1150 1999 1309 2001
rect 1111 1970 1113 1982
rect 1150 1970 1152 1999
rect 1345 1991 1347 2180
rect 1533 2176 1535 2180
rect 1533 2174 1754 2176
rect 1357 2169 1450 2171
rect 1448 2143 1450 2169
rect 1644 2167 1717 2169
rect 1379 2141 1382 2143
rect 1432 2141 1454 2143
rect 1474 2141 1477 2143
rect 1626 2133 1628 2139
rect 1556 2131 1559 2133
rect 1599 2131 1647 2133
rect 1687 2131 1690 2133
rect 1556 2092 1559 2094
rect 1599 2092 1647 2094
rect 1687 2092 1690 2094
rect 1448 2068 1450 2074
rect 1386 2066 1389 2068
rect 1429 2066 1477 2068
rect 1517 2066 1520 2068
rect 1635 2061 1637 2092
rect 1715 2064 1717 2167
rect 1752 2159 1754 2174
rect 1951 2202 1953 2211
rect 1990 2202 1992 2220
rect 1827 2159 1829 2163
rect 1752 2157 1829 2159
rect 1866 2083 1868 2163
rect 1951 2159 1953 2162
rect 1990 2159 1992 2162
rect 2026 2083 2028 2505
rect 2100 2390 2107 2392
rect 2066 2290 2068 2293
rect 2105 2290 2107 2390
rect 2066 2231 2068 2250
rect 2058 2229 2068 2231
rect 2066 2202 2068 2229
rect 2105 2202 2107 2250
rect 2066 2159 2068 2162
rect 2105 2159 2107 2162
rect 1866 2081 2028 2083
rect 1715 2062 1868 2064
rect 1630 2059 1637 2061
rect 1599 2033 1602 2035
rect 1622 2033 1644 2035
rect 1694 2033 1697 2035
rect 1386 2027 1389 2029
rect 1429 2027 1477 2029
rect 1517 2027 1520 2029
rect 1439 1996 1441 2027
rect 1452 2003 1461 2005
rect 1459 2001 1461 2003
rect 1626 2001 1628 2033
rect 1459 1999 1628 2001
rect 1439 1994 1446 1996
rect 1235 1989 1347 1991
rect 1204 1978 1206 1981
rect 1111 1882 1113 1930
rect 1150 1882 1152 1930
rect 1204 1906 1206 1928
rect 1204 1883 1206 1886
rect 1111 1817 1113 1842
rect 1150 1838 1152 1842
rect 1235 1817 1237 1989
rect 1827 1982 1829 1985
rect 1866 1982 1868 2062
rect 2138 2025 2140 2227
rect 2215 2034 2217 2524
rect 2250 2503 2252 2524
rect 2289 2541 2291 2551
rect 2289 2539 2334 2541
rect 2289 2503 2291 2539
rect 2250 2460 2252 2463
rect 2289 2460 2291 2463
rect 2320 2439 2322 2528
rect 2289 2437 2322 2439
rect 2250 2431 2252 2434
rect 2289 2431 2291 2437
rect 2332 2427 2334 2539
rect 2552 2432 2554 2435
rect 2591 2432 2593 2435
rect 2250 2343 2252 2391
rect 2289 2343 2291 2391
rect 2552 2363 2554 2392
rect 2546 2361 2554 2363
rect 2552 2344 2554 2361
rect 2591 2344 2593 2392
rect 2637 2363 2644 2365
rect 2250 2291 2252 2303
rect 2289 2300 2291 2303
rect 2552 2301 2554 2304
rect 2245 2289 2252 2291
rect 2245 2276 2247 2289
rect 2245 2274 2252 2276
rect 2332 2275 2334 2297
rect 2591 2292 2593 2304
rect 2591 2290 2633 2292
rect 2250 2261 2252 2274
rect 2289 2273 2334 2275
rect 2289 2261 2291 2273
rect 2361 2269 2363 2272
rect 2250 2173 2252 2221
rect 2289 2173 2291 2221
rect 2426 2262 2428 2265
rect 2465 2262 2467 2265
rect 2552 2262 2554 2265
rect 2591 2262 2593 2265
rect 2631 2257 2633 2290
rect 2361 2197 2363 2219
rect 2426 2204 2428 2222
rect 2421 2202 2428 2204
rect 2361 2174 2363 2177
rect 2426 2174 2428 2202
rect 2465 2174 2467 2222
rect 2552 2203 2554 2222
rect 2548 2201 2554 2203
rect 2552 2174 2554 2201
rect 2591 2188 2593 2222
rect 2642 2188 2644 2363
rect 2591 2186 2644 2188
rect 2591 2174 2593 2186
rect 2250 2130 2252 2133
rect 2289 2130 2291 2133
rect 2426 2131 2428 2134
rect 2465 2126 2467 2134
rect 2465 2124 2470 2126
rect 2250 2101 2252 2104
rect 2289 2101 2291 2104
rect 2468 2071 2470 2124
rect 2215 2032 2225 2034
rect 2250 2025 2252 2061
rect 2138 2023 2252 2025
rect 2250 2013 2252 2023
rect 2289 2051 2291 2061
rect 2508 2051 2510 2137
rect 2552 2131 2554 2134
rect 2591 2131 2593 2134
rect 2289 2049 2510 2051
rect 2289 2013 2291 2049
rect 1951 1983 1953 1986
rect 1990 1983 1992 1986
rect 2066 1983 2068 1986
rect 2105 1983 2107 1986
rect 1111 1815 1237 1817
rect 1243 1803 1245 1969
rect 1379 1968 1382 1970
rect 1432 1968 1454 1970
rect 1474 1968 1477 1970
rect 1147 1801 1245 1803
rect 1108 1773 1110 1777
rect 1147 1773 1149 1801
rect 1108 1716 1110 1733
rect 1075 1714 1110 1716
rect 1108 1685 1110 1714
rect 1147 1685 1149 1733
rect 1201 1729 1203 1732
rect 1201 1687 1203 1709
rect 1108 1632 1110 1645
rect 1147 1642 1149 1645
rect 1201 1634 1203 1637
rect 1102 1630 1110 1632
rect 1102 1576 1104 1630
rect 1270 1596 1272 1936
rect 1448 1913 1450 1968
rect 2250 1970 2252 1973
rect 2289 1970 2291 1973
rect 1827 1924 1829 1942
rect 1287 1911 1450 1913
rect 1770 1922 1829 1924
rect 1143 1594 1272 1596
rect 1102 1574 1106 1576
rect 1104 1572 1106 1574
rect 1143 1572 1145 1594
rect 1104 1484 1106 1532
rect 1143 1484 1145 1532
rect 1197 1528 1199 1531
rect 1197 1486 1199 1508
rect 1057 968 1059 1439
rect 1104 1432 1106 1444
rect 1143 1441 1145 1444
rect 1197 1433 1199 1436
rect 1098 1430 1106 1432
rect 1098 1402 1100 1430
rect 1318 1417 1320 1911
rect 1770 1875 1772 1922
rect 1827 1894 1829 1922
rect 1866 1934 1868 1942
rect 1951 1934 1953 1943
rect 1866 1932 1953 1934
rect 1866 1894 1868 1932
rect 1383 1873 1772 1875
rect 1143 1415 1320 1417
rect 1098 1400 1106 1402
rect 1104 1388 1106 1400
rect 1143 1388 1145 1415
rect 1197 1396 1199 1399
rect 1104 1300 1106 1348
rect 1143 1300 1145 1348
rect 1197 1324 1199 1346
rect 1197 1301 1199 1304
rect 1104 1258 1106 1260
rect 1102 1256 1106 1258
rect 1102 1203 1104 1256
rect 1143 1239 1145 1260
rect 1340 1227 1342 1713
rect 1143 1225 1342 1227
rect 1102 1201 1106 1203
rect 1104 1199 1106 1201
rect 1143 1199 1145 1225
rect 1104 1111 1106 1159
rect 1143 1111 1145 1159
rect 1197 1155 1199 1158
rect 1197 1113 1199 1135
rect 1104 1059 1106 1071
rect 1143 1067 1145 1071
rect 1197 1060 1199 1063
rect 1097 1057 1106 1059
rect 1097 1034 1099 1057
rect 1383 1034 1385 1873
rect 1827 1842 1829 1854
rect 1866 1851 1868 1854
rect 1827 1840 1849 1842
rect 1847 1757 1849 1840
rect 1910 1826 1912 1910
rect 1951 1895 1953 1932
rect 1990 1925 1992 1943
rect 1984 1923 1992 1925
rect 1990 1895 1992 1923
rect 2066 1916 2068 1943
rect 2058 1914 2068 1916
rect 2066 1895 2068 1914
rect 2105 1895 2107 1943
rect 2250 1931 2252 1934
rect 2289 1931 2291 1934
rect 1951 1852 1953 1855
rect 1990 1852 1992 1855
rect 2066 1852 2068 1855
rect 1910 1824 1992 1826
rect 1951 1813 1953 1816
rect 1990 1813 1992 1824
rect 1951 1757 1953 1773
rect 1847 1755 1953 1757
rect 1951 1725 1953 1755
rect 1990 1725 1992 1773
rect 2105 1755 2107 1855
rect 2100 1753 2107 1755
rect 1401 1702 1543 1704
rect 1541 1607 1543 1702
rect 1951 1682 1953 1685
rect 1990 1682 1992 1685
rect 1472 1605 1475 1607
rect 1525 1605 1547 1607
rect 1567 1605 1570 1607
rect 1541 1532 1543 1538
rect 1479 1530 1482 1532
rect 1522 1530 1570 1532
rect 1610 1530 1613 1532
rect 1479 1491 1482 1493
rect 1522 1491 1570 1493
rect 1610 1491 1613 1493
rect 1532 1460 1534 1491
rect 1545 1468 1555 1470
rect 1532 1458 1539 1460
rect 1553 1458 1555 1468
rect 1553 1456 1725 1458
rect 1723 1437 1725 1456
rect 1696 1435 1699 1437
rect 1719 1435 1741 1437
rect 1791 1435 1794 1437
rect 1472 1432 1475 1434
rect 1525 1432 1547 1434
rect 1567 1432 1570 1434
rect 1541 1418 1543 1432
rect 1431 1416 1543 1418
rect 1754 1401 1824 1403
rect 1453 1398 1548 1400
rect 1546 1372 1548 1398
rect 1476 1370 1479 1372
rect 1529 1370 1551 1372
rect 1571 1370 1574 1372
rect 1723 1362 1725 1368
rect 1653 1360 1656 1362
rect 1696 1360 1744 1362
rect 1784 1360 1787 1362
rect 1653 1321 1656 1323
rect 1696 1321 1744 1323
rect 1784 1321 1787 1323
rect 1545 1297 1547 1303
rect 1483 1295 1486 1297
rect 1526 1295 1574 1297
rect 1614 1295 1617 1297
rect 1732 1290 1734 1321
rect 1727 1288 1734 1290
rect 1696 1262 1699 1264
rect 1719 1262 1741 1264
rect 1791 1262 1794 1264
rect 1483 1256 1486 1258
rect 1526 1256 1574 1258
rect 1614 1256 1617 1258
rect 1536 1225 1538 1256
rect 1549 1232 1558 1234
rect 1556 1230 1558 1232
rect 1723 1230 1725 1262
rect 1556 1228 1725 1230
rect 1536 1223 1543 1225
rect 1822 1203 1824 1401
rect 2140 1365 2142 1911
rect 2250 1866 2252 1891
rect 2215 1864 2252 1866
rect 2215 1374 2217 1864
rect 2250 1843 2252 1864
rect 2289 1881 2291 1891
rect 2289 1879 2334 1881
rect 2289 1843 2291 1879
rect 2250 1800 2252 1803
rect 2289 1800 2291 1803
rect 2320 1779 2322 1868
rect 2289 1777 2322 1779
rect 2250 1771 2252 1774
rect 2289 1771 2291 1777
rect 2332 1767 2334 1879
rect 2552 1772 2554 1775
rect 2591 1772 2593 1775
rect 2250 1683 2252 1731
rect 2289 1683 2291 1731
rect 2552 1703 2554 1732
rect 2546 1701 2554 1703
rect 2552 1684 2554 1701
rect 2591 1684 2593 1732
rect 2637 1703 2644 1705
rect 2250 1631 2252 1643
rect 2289 1640 2291 1643
rect 2552 1641 2554 1644
rect 2245 1629 2252 1631
rect 2245 1616 2247 1629
rect 2245 1614 2252 1616
rect 2332 1615 2334 1637
rect 2591 1632 2593 1644
rect 2591 1630 2633 1632
rect 2250 1601 2252 1614
rect 2289 1613 2334 1615
rect 2289 1601 2291 1613
rect 2361 1609 2363 1612
rect 2250 1513 2252 1561
rect 2289 1513 2291 1561
rect 2426 1602 2428 1605
rect 2465 1602 2467 1605
rect 2552 1602 2554 1605
rect 2591 1602 2593 1605
rect 2631 1597 2633 1630
rect 2361 1537 2363 1559
rect 2426 1544 2428 1562
rect 2421 1542 2428 1544
rect 2361 1514 2363 1517
rect 2426 1514 2428 1542
rect 2465 1514 2467 1562
rect 2552 1543 2554 1562
rect 2548 1541 2554 1543
rect 2552 1514 2554 1541
rect 2591 1528 2593 1562
rect 2642 1528 2644 1703
rect 2591 1526 2644 1528
rect 2591 1514 2593 1526
rect 2250 1470 2252 1473
rect 2289 1470 2291 1473
rect 2426 1471 2428 1474
rect 2465 1466 2467 1474
rect 2465 1464 2470 1466
rect 2250 1441 2252 1444
rect 2289 1441 2291 1444
rect 2468 1411 2470 1464
rect 2215 1372 2225 1374
rect 2250 1365 2252 1401
rect 2140 1363 2252 1365
rect 2250 1353 2252 1363
rect 2289 1391 2291 1401
rect 2508 1391 2510 1477
rect 2552 1471 2554 1474
rect 2591 1471 2593 1474
rect 2289 1389 2510 1391
rect 2289 1353 2291 1389
rect 2250 1310 2252 1313
rect 2289 1310 2291 1313
rect 2250 1271 2252 1274
rect 2289 1271 2291 1274
rect 2250 1206 2252 1231
rect 1714 1201 1824 1203
rect 2215 1204 2252 1206
rect 1476 1197 1479 1199
rect 1529 1197 1551 1199
rect 1571 1197 1574 1199
rect 1545 1130 1547 1197
rect 1714 1175 1716 1201
rect 1687 1173 1690 1175
rect 1710 1173 1732 1175
rect 1782 1173 1785 1175
rect 1729 1145 1814 1147
rect 1424 1128 1547 1130
rect 1714 1100 1716 1106
rect 1644 1098 1647 1100
rect 1687 1098 1735 1100
rect 1775 1098 1778 1100
rect 1644 1059 1647 1061
rect 1687 1059 1735 1061
rect 1775 1059 1778 1061
rect 1097 1032 1385 1034
rect 1723 1028 1725 1059
rect 1718 1026 1725 1028
rect 1687 1000 1690 1002
rect 1710 1000 1732 1002
rect 1782 1000 1785 1002
rect 1714 968 1716 1000
rect 1057 966 1716 968
rect 1812 705 1814 1145
rect 2215 714 2217 1204
rect 2250 1183 2252 1204
rect 2289 1221 2291 1231
rect 2289 1219 2334 1221
rect 2289 1183 2291 1219
rect 2250 1140 2252 1143
rect 2289 1140 2291 1143
rect 2320 1119 2322 1208
rect 2289 1117 2322 1119
rect 2250 1111 2252 1114
rect 2289 1111 2291 1117
rect 2332 1107 2334 1219
rect 2552 1112 2554 1115
rect 2591 1112 2593 1115
rect 2250 1023 2252 1071
rect 2289 1023 2291 1071
rect 2552 1043 2554 1072
rect 2546 1041 2554 1043
rect 2552 1024 2554 1041
rect 2591 1024 2593 1072
rect 2637 1043 2644 1045
rect 2250 971 2252 983
rect 2289 980 2291 983
rect 2552 981 2554 984
rect 2245 969 2252 971
rect 2245 956 2247 969
rect 2245 954 2252 956
rect 2332 955 2334 977
rect 2591 972 2593 984
rect 2591 970 2633 972
rect 2250 941 2252 954
rect 2289 953 2334 955
rect 2289 941 2291 953
rect 2361 949 2363 952
rect 2250 853 2252 901
rect 2289 853 2291 901
rect 2426 942 2428 945
rect 2465 942 2467 945
rect 2552 942 2554 945
rect 2591 942 2593 945
rect 2631 937 2633 970
rect 2361 877 2363 899
rect 2426 884 2428 902
rect 2421 882 2428 884
rect 2361 854 2363 857
rect 2426 854 2428 882
rect 2465 854 2467 902
rect 2552 883 2554 902
rect 2548 881 2554 883
rect 2552 854 2554 881
rect 2591 868 2593 902
rect 2642 868 2644 1043
rect 2591 866 2644 868
rect 2591 854 2593 866
rect 2250 810 2252 813
rect 2289 810 2291 813
rect 2426 811 2428 814
rect 2465 806 2467 814
rect 2465 804 2470 806
rect 2250 781 2252 784
rect 2289 781 2291 784
rect 2468 751 2470 804
rect 2215 712 2225 714
rect 2250 705 2252 741
rect 1812 703 2252 705
rect 2250 693 2252 703
rect 2289 731 2291 741
rect 2508 731 2510 817
rect 2552 811 2554 814
rect 2591 811 2593 814
rect 2289 729 2510 731
rect 2289 693 2291 729
rect 2250 650 2252 653
rect 2289 650 2291 653
rect 436 156 959 158
rect 100 151 188 153
rect 252 109 254 113
rect 182 107 185 109
rect 225 107 273 109
rect 313 107 316 109
rect 412 109 414 115
rect 352 107 355 109
rect 395 107 443 109
rect 483 107 486 109
rect 182 68 185 70
rect 225 68 273 70
rect 313 68 316 70
rect 341 68 355 70
rect 395 68 443 70
rect 483 68 486 70
rect 237 19 239 68
rect 341 30 343 68
rect 308 28 343 30
rect 414 19 416 24
rect 237 17 416 19
<< polycontact >>
rect 80 4261 87 4267
rect 579 4167 586 4174
rect 348 4156 355 4162
rect 473 4156 478 4162
rect 251 4131 256 4136
rect 251 4071 256 4075
rect 116 4018 122 4026
rect 430 3985 436 3991
rect 188 3980 192 3985
rect 250 3944 257 3949
rect 410 3946 417 3951
rect 303 3857 308 3863
rect 411 3855 418 3860
rect 430 3507 436 3513
rect 1163 3623 1168 3628
rect 1177 3591 1181 3596
rect 1163 3554 1168 3558
rect 80 3304 87 3310
rect 1163 3473 1168 3477
rect 1264 3424 1268 3428
rect 1066 3378 1071 3386
rect 1164 3290 1169 3295
rect 579 3210 586 3217
rect 348 3199 355 3205
rect 473 3199 478 3205
rect 251 3174 256 3179
rect 251 3114 256 3118
rect 116 3061 122 3069
rect 430 3028 436 3034
rect 1908 3356 1915 3361
rect 1980 3344 1984 3350
rect 2095 3514 2100 3521
rect 2053 3353 2058 3360
rect 2134 3353 2140 3360
rect 2318 3848 2325 3855
rect 2330 3742 2336 3747
rect 2541 3679 2546 3686
rect 2632 3680 2637 3687
rect 2330 3617 2336 3624
rect 2629 3572 2635 3577
rect 2356 3520 2361 3525
rect 2417 3520 2421 3525
rect 2543 3519 2548 3526
rect 2507 3457 2512 3461
rect 2466 3385 2474 3391
rect 2225 3349 2231 3356
rect 188 3023 192 3028
rect 838 3156 845 3161
rect 910 3167 914 3173
rect 983 3157 988 3164
rect 1066 3157 1071 3165
rect 1164 3162 1169 3167
rect 829 3043 835 3049
rect 250 2987 257 2992
rect 410 2989 417 2994
rect 303 2900 308 2906
rect 411 2898 418 2903
rect 80 2825 87 2831
rect 579 2731 586 2738
rect 348 2720 355 2726
rect 473 2720 478 2726
rect 251 2695 256 2700
rect 251 2635 256 2639
rect 116 2582 122 2590
rect 430 2549 436 2555
rect 792 2832 798 2837
rect 779 2774 784 2779
rect 1025 2996 1030 3003
rect 1173 3069 1178 3074
rect 1908 3036 1915 3041
rect 1285 3000 1290 3005
rect 1980 3047 1984 3053
rect 2053 3037 2058 3044
rect 2138 3037 2144 3044
rect 1174 2864 1179 2869
rect 2095 2876 2100 2883
rect 1225 2825 1229 2830
rect 1174 2783 1179 2788
rect 188 2544 192 2549
rect 250 2508 257 2513
rect 410 2510 417 2515
rect 303 2421 308 2427
rect 411 2419 418 2424
rect 80 2346 87 2352
rect 579 2252 586 2259
rect 348 2241 355 2247
rect 473 2241 478 2247
rect 251 2216 256 2221
rect 251 2156 256 2160
rect 116 2103 122 2111
rect 430 2070 436 2076
rect 1174 2714 1179 2718
rect 779 2638 784 2643
rect 1174 2633 1179 2637
rect 1174 2603 1179 2608
rect 792 2580 798 2585
rect 1148 2567 1153 2571
rect 1025 2414 1030 2421
rect 829 2368 835 2374
rect 838 2256 845 2261
rect 910 2244 914 2250
rect 983 2253 988 2260
rect 188 2065 192 2070
rect 250 2029 257 2034
rect 410 2031 417 2036
rect 303 1942 308 1948
rect 411 1940 418 1945
rect 80 1867 87 1873
rect 579 1773 586 1780
rect 348 1762 355 1768
rect 473 1762 478 1768
rect 1066 2252 1071 2260
rect 1199 2255 1204 2260
rect 1379 2733 1384 2738
rect 2318 3188 2325 3195
rect 2330 3082 2336 3087
rect 2541 3019 2546 3026
rect 2632 3020 2637 3027
rect 2330 2957 2336 2964
rect 2629 2912 2635 2917
rect 2356 2860 2361 2865
rect 2417 2860 2421 2865
rect 2543 2859 2548 2866
rect 2507 2797 2512 2801
rect 2466 2725 2474 2731
rect 2225 2689 2231 2696
rect 1379 2664 1384 2668
rect 1378 2592 1385 2597
rect 1379 2583 1384 2587
rect 1379 2553 1384 2558
rect 1305 2522 1311 2526
rect 251 1737 256 1742
rect 251 1677 256 1681
rect 116 1624 122 1632
rect 430 1591 436 1597
rect 1199 2084 1204 2089
rect 838 2030 845 2035
rect 910 2041 914 2047
rect 983 2031 988 2038
rect 1066 2031 1071 2039
rect 829 1917 835 1923
rect 188 1586 192 1591
rect 250 1550 257 1555
rect 410 1552 417 1557
rect 303 1463 308 1469
rect 411 1461 418 1466
rect 80 1388 87 1394
rect 579 1294 586 1301
rect 348 1283 355 1289
rect 473 1283 478 1289
rect 251 1258 256 1263
rect 251 1198 256 1202
rect 116 1145 122 1153
rect 430 1112 436 1118
rect 792 1706 798 1711
rect 779 1648 784 1653
rect 188 1107 192 1112
rect 250 1071 257 1076
rect 410 1073 417 1078
rect 303 984 308 990
rect 411 982 418 987
rect 80 909 87 915
rect 579 815 586 822
rect 348 804 355 810
rect 473 804 478 810
rect 251 779 256 784
rect 251 719 256 723
rect 116 666 122 674
rect 430 633 436 639
rect 188 628 192 633
rect 250 592 257 597
rect 410 594 417 599
rect 303 505 308 511
rect 411 503 418 508
rect 80 430 87 436
rect 579 336 586 343
rect 348 325 355 331
rect 473 325 478 331
rect 251 300 256 305
rect 251 240 256 244
rect 116 187 122 195
rect 430 154 436 160
rect 1025 1870 1030 1877
rect 1318 2404 1322 2410
rect 1442 2309 1447 2313
rect 1441 2238 1448 2243
rect 1442 2228 1447 2232
rect 1908 2230 1915 2235
rect 1980 2218 1984 2224
rect 1313 2175 1317 2179
rect 1352 2168 1357 2172
rect 1640 2165 1644 2170
rect 1625 2139 1630 2143
rect 1446 2074 1451 2078
rect 1625 2058 1630 2062
rect 2095 2388 2100 2395
rect 2053 2227 2058 2234
rect 2136 2227 2142 2234
rect 1445 2001 1452 2007
rect 1446 1993 1451 1997
rect 1199 1909 1204 1914
rect 2318 2528 2325 2535
rect 2330 2422 2336 2427
rect 2541 2359 2546 2366
rect 2632 2360 2637 2367
rect 2330 2297 2336 2304
rect 2629 2252 2635 2257
rect 2356 2200 2361 2205
rect 2417 2200 2421 2205
rect 2543 2199 2548 2206
rect 2507 2137 2512 2141
rect 2466 2065 2474 2071
rect 2225 2029 2231 2036
rect 1241 1969 1246 1973
rect 1268 1936 1273 1941
rect 1196 1701 1201 1706
rect 1283 1909 1287 1914
rect 1192 1500 1197 1505
rect 1056 1439 1061 1443
rect 1908 1910 1915 1915
rect 1339 1713 1343 1717
rect 1192 1327 1197 1332
rect 1192 1127 1197 1132
rect 1980 1921 1984 1927
rect 2053 1911 2058 1918
rect 2138 1911 2143 1918
rect 2095 1750 2100 1757
rect 1395 1701 1401 1706
rect 1539 1538 1544 1542
rect 1538 1467 1545 1472
rect 1539 1457 1544 1461
rect 1425 1415 1431 1420
rect 1448 1397 1453 1401
rect 1750 1400 1754 1404
rect 1722 1368 1727 1372
rect 1543 1303 1548 1307
rect 1722 1287 1727 1291
rect 1542 1230 1549 1236
rect 1543 1222 1548 1226
rect 2318 1868 2325 1875
rect 2330 1762 2336 1767
rect 2541 1699 2546 1706
rect 2632 1700 2637 1707
rect 2330 1637 2336 1644
rect 2629 1592 2635 1597
rect 2356 1540 2361 1545
rect 2417 1540 2421 1545
rect 2543 1539 2548 1546
rect 2507 1477 2512 1481
rect 2466 1405 2474 1411
rect 2225 1369 2231 1376
rect 1419 1127 1424 1132
rect 1725 1144 1729 1148
rect 1713 1106 1718 1110
rect 1713 1025 1718 1029
rect 2318 1208 2325 1215
rect 2330 1102 2336 1107
rect 2541 1039 2546 1046
rect 2632 1040 2637 1047
rect 2330 977 2336 984
rect 2629 932 2635 937
rect 2356 880 2361 885
rect 2417 880 2421 885
rect 2543 879 2548 886
rect 2507 817 2512 821
rect 2466 745 2474 751
rect 2225 709 2231 716
rect 188 149 192 154
rect 250 113 257 118
rect 410 115 417 120
rect 303 26 308 32
rect 411 24 418 29
<< metal1 >>
rect 0 4309 727 4315
rect 0 4259 6 4309
rect 165 4284 501 4290
rect 0 4252 26 4259
rect 0 4243 6 4252
rect 0 4192 6 4235
rect 80 4225 87 4261
rect 165 4259 171 4284
rect 495 4259 501 4284
rect 660 4259 666 4309
rect 150 4252 186 4259
rect 310 4252 356 4259
rect 480 4252 516 4259
rect 640 4252 666 4259
rect 64 4218 87 4225
rect 80 4193 87 4218
rect 165 4231 171 4252
rect 330 4243 336 4252
rect 0 4185 26 4192
rect 80 4186 112 4193
rect 0 3836 6 4185
rect 80 4026 87 4186
rect 165 4151 171 4223
rect 249 4218 272 4225
rect 249 4193 256 4218
rect 224 4186 256 4193
rect 330 4192 336 4235
rect 495 4231 501 4252
rect 394 4218 417 4225
rect 410 4193 417 4218
rect 660 4243 666 4252
rect 165 4146 224 4151
rect 165 4083 171 4146
rect 219 4136 224 4146
rect 251 4136 256 4186
rect 310 4185 356 4192
rect 410 4186 442 4193
rect 332 4136 337 4185
rect 410 4162 417 4186
rect 355 4156 473 4162
rect 219 4132 228 4136
rect 219 4102 224 4132
rect 320 4132 337 4136
rect 248 4124 270 4128
rect 165 4082 187 4083
rect 166 4076 187 4082
rect 166 4055 172 4076
rect 251 4075 256 4124
rect 332 4083 337 4132
rect 311 4076 337 4083
rect 331 4067 337 4076
rect 80 4018 116 4026
rect 166 3957 172 4047
rect 250 4042 273 4049
rect 250 4017 257 4042
rect 225 4010 257 4017
rect 331 4016 337 4059
rect 250 3985 257 4010
rect 311 4009 337 4016
rect 192 3980 257 3985
rect 166 3950 187 3957
rect 166 3929 172 3950
rect 250 3949 257 3980
rect 331 3957 337 4009
rect 311 3950 357 3957
rect 410 3951 417 4156
rect 331 3941 337 3950
rect 166 3883 172 3921
rect 250 3916 273 3923
rect 250 3891 257 3916
rect 225 3884 257 3891
rect 331 3890 337 3933
rect 430 3923 436 3985
rect 495 3957 501 4223
rect 579 4218 602 4225
rect 579 4193 586 4218
rect 554 4186 586 4193
rect 660 4192 666 4235
rect 579 4174 586 4186
rect 640 4185 666 4192
rect 481 3950 502 3957
rect 395 3916 436 3923
rect 496 3929 502 3950
rect 411 3891 418 3916
rect 250 3863 257 3884
rect 311 3883 357 3890
rect 411 3884 443 3891
rect 496 3888 502 3921
rect 250 3857 303 3863
rect 331 3836 337 3883
rect 411 3860 418 3884
rect 496 3883 676 3888
rect 0 3831 337 3836
rect 430 3445 436 3507
rect 417 3438 436 3445
rect 671 3410 676 3883
rect 721 3837 727 4309
rect 2177 3929 2249 3935
rect 2257 3929 2307 3935
rect 2177 3837 2183 3929
rect 2233 3909 2240 3929
rect 2300 3909 2307 3929
rect 2267 3855 2274 3871
rect 2267 3848 2318 3855
rect 698 3832 2183 3837
rect 698 3781 703 3832
rect 779 3816 1168 3822
rect 779 3795 784 3816
rect 1163 3645 1168 3816
rect 1078 3598 1083 3633
rect 1131 3628 1136 3643
rect 1163 3639 1343 3645
rect 1163 3628 1168 3639
rect 1244 3628 1249 3635
rect 1131 3624 1140 3628
rect 1131 3598 1136 3624
rect 1232 3624 1249 3628
rect 1160 3616 1182 3620
rect 1078 3594 1136 3598
rect 1078 3565 1083 3594
rect 1078 3558 1099 3565
rect 1163 3558 1168 3616
rect 1078 3537 1084 3558
rect 1171 3591 1177 3596
rect 1171 3531 1176 3591
rect 1244 3565 1249 3624
rect 1223 3558 1249 3565
rect 1243 3549 1249 3558
rect 1078 3491 1084 3529
rect 1162 3524 1185 3531
rect 1162 3499 1169 3524
rect 1137 3492 1169 3499
rect 1243 3498 1249 3541
rect 1223 3491 1249 3498
rect 502 3405 676 3410
rect 0 3352 666 3358
rect 0 3302 6 3352
rect 165 3327 501 3333
rect 0 3295 26 3302
rect 0 3286 6 3295
rect 0 3235 6 3278
rect 80 3268 87 3304
rect 165 3302 171 3327
rect 495 3302 501 3327
rect 660 3302 666 3352
rect 150 3295 186 3302
rect 310 3295 356 3302
rect 480 3295 516 3302
rect 640 3295 666 3302
rect 64 3261 87 3268
rect 80 3236 87 3261
rect 165 3274 171 3295
rect 330 3286 336 3295
rect 0 3228 26 3235
rect 80 3229 112 3236
rect 0 2879 6 3228
rect 80 3069 87 3229
rect 165 3194 171 3266
rect 249 3261 272 3268
rect 249 3236 256 3261
rect 224 3229 256 3236
rect 330 3235 336 3278
rect 495 3274 501 3295
rect 394 3261 417 3268
rect 410 3236 417 3261
rect 660 3286 666 3295
rect 165 3189 224 3194
rect 165 3126 171 3189
rect 219 3179 224 3189
rect 251 3179 256 3229
rect 310 3228 356 3235
rect 410 3229 442 3236
rect 332 3179 337 3228
rect 410 3205 417 3229
rect 355 3199 473 3205
rect 219 3175 228 3179
rect 219 3145 224 3175
rect 320 3175 337 3179
rect 248 3167 270 3171
rect 165 3125 187 3126
rect 166 3119 187 3125
rect 166 3098 172 3119
rect 251 3118 256 3167
rect 332 3126 337 3175
rect 311 3119 337 3126
rect 331 3110 337 3119
rect 80 3061 116 3069
rect 166 3000 172 3090
rect 250 3085 273 3092
rect 250 3060 257 3085
rect 225 3053 257 3060
rect 331 3059 337 3102
rect 250 3028 257 3053
rect 311 3052 337 3059
rect 192 3023 257 3028
rect 166 2993 187 3000
rect 166 2972 172 2993
rect 250 2992 257 3023
rect 331 3000 337 3052
rect 311 2993 357 3000
rect 410 2994 417 3199
rect 331 2984 337 2993
rect 166 2926 172 2964
rect 250 2959 273 2966
rect 250 2934 257 2959
rect 225 2927 257 2934
rect 331 2933 337 2976
rect 430 2966 436 3028
rect 495 3000 501 3266
rect 579 3261 602 3268
rect 579 3236 586 3261
rect 554 3229 586 3236
rect 660 3235 666 3278
rect 579 3217 586 3229
rect 640 3228 666 3235
rect 481 2993 502 3000
rect 395 2959 436 2966
rect 496 2972 502 2993
rect 671 2985 676 3405
rect 699 3082 705 3462
rect 1078 3451 1083 3491
rect 1244 3484 1249 3491
rect 1244 3477 1319 3484
rect 1163 3455 1168 3473
rect 1131 3451 1136 3453
rect 1160 3451 1182 3455
rect 1078 3447 1136 3451
rect 1244 3447 1249 3477
rect 1078 3445 1083 3447
rect 1131 3443 1140 3447
rect 1232 3443 1249 3447
rect 1131 3441 1136 3443
rect 1244 3400 1249 3443
rect 1268 3424 1281 3428
rect 1078 3393 1099 3400
rect 1223 3393 1249 3400
rect 1059 3378 1066 3386
rect 1078 3372 1084 3393
rect 1243 3384 1249 3393
rect 1078 3310 1084 3364
rect 1162 3359 1185 3366
rect 1162 3334 1169 3359
rect 1137 3327 1169 3334
rect 1243 3333 1249 3376
rect 1078 3305 1137 3310
rect 1132 3295 1137 3305
rect 1164 3295 1169 3327
rect 1223 3327 1249 3333
rect 1223 3326 1250 3327
rect 1245 3295 1250 3326
rect 1132 3291 1141 3295
rect 1132 3248 1137 3291
rect 1233 3291 1250 3295
rect 1161 3283 1183 3287
rect 864 3247 892 3248
rect 740 3241 768 3247
rect 776 3242 892 3247
rect 900 3242 1007 3248
rect 1015 3242 1137 3248
rect 1164 3256 1169 3283
rect 1245 3277 1250 3291
rect 1276 3256 1281 3424
rect 1164 3252 1281 3256
rect 776 3241 871 3242
rect 740 3226 747 3241
rect 864 3227 871 3241
rect 979 3227 986 3242
rect 806 3173 813 3188
rect 806 3167 910 3173
rect 806 3163 813 3167
rect 774 3156 813 3163
rect 838 3161 845 3167
rect 930 3164 937 3189
rect 1045 3165 1052 3189
rect 1087 3179 1092 3242
rect 1087 3172 1108 3179
rect 1045 3164 1066 3165
rect 898 3157 983 3164
rect 1013 3157 1066 3164
rect 774 3140 781 3156
rect 898 3141 905 3157
rect 1013 3141 1020 3157
rect 1087 3151 1093 3172
rect 1164 3167 1169 3252
rect 1312 3179 1319 3477
rect 1232 3172 1319 3179
rect 1252 3163 1258 3172
rect 740 3082 747 3102
rect 807 3083 814 3102
rect 864 3083 871 3103
rect 931 3083 938 3103
rect 979 3083 986 3103
rect 1046 3083 1053 3103
rect 807 3082 880 3083
rect 699 3076 756 3082
rect 764 3077 880 3082
rect 888 3077 995 3083
rect 1003 3077 1053 3083
rect 1087 3089 1093 3143
rect 1171 3138 1194 3145
rect 1171 3113 1178 3138
rect 1146 3106 1178 3113
rect 1252 3112 1258 3155
rect 1087 3084 1146 3089
rect 764 3076 871 3077
rect 671 2980 688 2985
rect 411 2934 418 2959
rect 250 2906 257 2927
rect 311 2926 357 2933
rect 411 2927 443 2934
rect 496 2931 502 2964
rect 684 2931 688 2980
rect 250 2900 303 2906
rect 331 2879 337 2926
rect 411 2903 418 2927
rect 496 2926 688 2931
rect 0 2873 666 2879
rect 0 2823 6 2873
rect 165 2848 501 2854
rect 0 2816 26 2823
rect 0 2807 6 2816
rect 0 2756 6 2799
rect 80 2789 87 2825
rect 165 2823 171 2848
rect 495 2823 501 2848
rect 660 2823 666 2873
rect 150 2816 186 2823
rect 310 2816 356 2823
rect 480 2816 516 2823
rect 640 2816 666 2823
rect 64 2782 87 2789
rect 80 2757 87 2782
rect 165 2795 171 2816
rect 330 2807 336 2816
rect 0 2749 26 2756
rect 80 2750 112 2757
rect 0 2400 6 2749
rect 80 2590 87 2750
rect 165 2715 171 2787
rect 249 2782 272 2789
rect 249 2757 256 2782
rect 224 2750 256 2757
rect 330 2756 336 2799
rect 495 2795 501 2816
rect 394 2782 417 2789
rect 410 2757 417 2782
rect 660 2807 666 2816
rect 165 2710 224 2715
rect 165 2647 171 2710
rect 219 2700 224 2710
rect 251 2700 256 2750
rect 310 2749 356 2756
rect 410 2750 442 2757
rect 332 2700 337 2749
rect 410 2726 417 2750
rect 355 2720 473 2726
rect 219 2696 228 2700
rect 219 2666 224 2696
rect 320 2696 337 2700
rect 248 2688 270 2692
rect 165 2646 187 2647
rect 166 2640 187 2646
rect 166 2619 172 2640
rect 251 2639 256 2688
rect 332 2647 337 2696
rect 311 2640 337 2647
rect 331 2631 337 2640
rect 80 2582 116 2590
rect 166 2521 172 2611
rect 250 2606 273 2613
rect 250 2581 257 2606
rect 225 2574 257 2581
rect 331 2580 337 2623
rect 250 2549 257 2574
rect 311 2573 337 2580
rect 192 2544 257 2549
rect 166 2514 187 2521
rect 166 2493 172 2514
rect 250 2513 257 2544
rect 331 2521 337 2573
rect 311 2514 357 2521
rect 410 2515 417 2720
rect 331 2505 337 2514
rect 166 2447 172 2485
rect 250 2480 273 2487
rect 250 2455 257 2480
rect 225 2448 257 2455
rect 331 2454 337 2497
rect 430 2487 436 2549
rect 495 2521 501 2787
rect 579 2782 602 2789
rect 579 2757 586 2782
rect 554 2750 586 2757
rect 660 2756 666 2799
rect 579 2738 586 2750
rect 640 2749 666 2756
rect 481 2514 502 2521
rect 395 2480 436 2487
rect 496 2493 502 2514
rect 411 2455 418 2480
rect 250 2427 257 2448
rect 311 2447 357 2454
rect 411 2448 443 2455
rect 496 2452 502 2485
rect 684 2452 688 2926
rect 699 2884 705 3076
rect 864 3057 871 3076
rect 931 3057 938 3077
rect 829 2970 835 3043
rect 1087 3051 1093 3084
rect 1141 3074 1146 3084
rect 1173 3074 1178 3106
rect 1232 3106 1258 3112
rect 1232 3105 1259 3106
rect 1254 3074 1259 3105
rect 1141 3070 1150 3074
rect 1141 3063 1146 3070
rect 1242 3070 1259 3074
rect 1170 3062 1192 3066
rect 1046 3045 1093 3051
rect 898 3003 905 3019
rect 898 2996 1025 3003
rect 930 2971 937 2996
rect 802 2966 835 2970
rect 699 2877 725 2884
rect 699 2868 705 2877
rect 699 2817 705 2860
rect 802 2858 806 2966
rect 864 2918 871 2933
rect 1046 2918 1052 3045
rect 1173 3035 1178 3062
rect 864 2912 892 2918
rect 900 2912 1052 2918
rect 1063 3031 1178 3035
rect 864 2884 870 2912
rect 849 2877 870 2884
rect 792 2854 806 2858
rect 864 2856 870 2877
rect 763 2843 786 2850
rect 779 2818 786 2843
rect 792 2837 798 2854
rect 699 2811 725 2817
rect 698 2810 725 2811
rect 779 2811 811 2818
rect 698 2779 703 2810
rect 779 2779 784 2811
rect 864 2794 870 2848
rect 811 2789 870 2794
rect 811 2779 816 2789
rect 698 2775 715 2779
rect 698 2711 703 2775
rect 807 2775 816 2779
rect 765 2767 787 2771
rect 779 2727 784 2767
rect 811 2765 816 2775
rect 779 2721 1052 2727
rect 698 2706 1036 2711
rect 698 2642 703 2706
rect 779 2675 1017 2681
rect 779 2650 784 2675
rect 765 2646 787 2650
rect 698 2638 715 2642
rect 811 2642 816 2655
rect 807 2638 816 2642
rect 698 2607 703 2638
rect 698 2606 725 2607
rect 250 2421 303 2427
rect 331 2400 337 2447
rect 411 2424 418 2448
rect 496 2447 688 2452
rect 0 2394 666 2400
rect 0 2344 6 2394
rect 165 2369 501 2375
rect 0 2337 26 2344
rect 0 2328 6 2337
rect 0 2277 6 2320
rect 80 2310 87 2346
rect 165 2344 171 2369
rect 495 2344 501 2369
rect 660 2344 666 2394
rect 150 2337 186 2344
rect 310 2337 356 2344
rect 480 2337 516 2344
rect 640 2337 666 2344
rect 64 2303 87 2310
rect 80 2278 87 2303
rect 165 2316 171 2337
rect 330 2328 336 2337
rect 0 2270 26 2277
rect 80 2271 112 2278
rect 0 1921 6 2270
rect 80 2111 87 2271
rect 165 2236 171 2308
rect 249 2303 272 2310
rect 249 2278 256 2303
rect 224 2271 256 2278
rect 330 2277 336 2320
rect 495 2316 501 2337
rect 394 2303 417 2310
rect 410 2278 417 2303
rect 660 2328 666 2337
rect 165 2231 224 2236
rect 165 2168 171 2231
rect 219 2221 224 2231
rect 251 2221 256 2271
rect 310 2270 356 2277
rect 410 2271 442 2278
rect 332 2221 337 2270
rect 410 2247 417 2271
rect 355 2241 473 2247
rect 219 2217 228 2221
rect 219 2187 224 2217
rect 320 2217 337 2221
rect 248 2209 270 2213
rect 165 2167 187 2168
rect 166 2161 187 2167
rect 166 2140 172 2161
rect 251 2160 256 2209
rect 332 2168 337 2217
rect 311 2161 337 2168
rect 331 2152 337 2161
rect 80 2103 116 2111
rect 166 2042 172 2132
rect 250 2127 273 2134
rect 250 2102 257 2127
rect 225 2095 257 2102
rect 331 2101 337 2144
rect 250 2070 257 2095
rect 311 2094 337 2101
rect 192 2065 257 2070
rect 166 2035 187 2042
rect 166 2014 172 2035
rect 250 2034 257 2065
rect 331 2042 337 2094
rect 311 2035 357 2042
rect 410 2036 417 2241
rect 331 2026 337 2035
rect 166 1968 172 2006
rect 250 2001 273 2008
rect 250 1976 257 2001
rect 225 1969 257 1976
rect 331 1975 337 2018
rect 430 2008 436 2070
rect 495 2042 501 2308
rect 579 2303 602 2310
rect 579 2278 586 2303
rect 554 2271 586 2278
rect 660 2277 666 2320
rect 579 2259 586 2271
rect 640 2270 666 2277
rect 481 2035 502 2042
rect 395 2001 436 2008
rect 496 2014 502 2035
rect 411 1976 418 2001
rect 250 1948 257 1969
rect 311 1968 357 1975
rect 411 1969 443 1976
rect 496 1973 502 2006
rect 684 1973 688 2447
rect 250 1942 303 1948
rect 331 1921 337 1968
rect 411 1945 418 1969
rect 496 1968 688 1973
rect 0 1915 666 1921
rect 0 1865 6 1915
rect 165 1890 501 1896
rect 0 1858 26 1865
rect 0 1849 6 1858
rect 0 1798 6 1841
rect 80 1831 87 1867
rect 165 1865 171 1890
rect 495 1865 501 1890
rect 660 1865 666 1915
rect 150 1858 186 1865
rect 310 1858 356 1865
rect 480 1858 516 1865
rect 640 1858 666 1865
rect 64 1824 87 1831
rect 80 1799 87 1824
rect 165 1837 171 1858
rect 330 1849 336 1858
rect 0 1791 26 1798
rect 80 1792 112 1799
rect 0 1442 6 1791
rect 80 1632 87 1792
rect 165 1757 171 1829
rect 249 1824 272 1831
rect 249 1799 256 1824
rect 224 1792 256 1799
rect 330 1798 336 1841
rect 495 1837 501 1858
rect 394 1824 417 1831
rect 410 1799 417 1824
rect 660 1849 666 1858
rect 165 1752 224 1757
rect 165 1689 171 1752
rect 219 1742 224 1752
rect 251 1742 256 1792
rect 310 1791 356 1798
rect 410 1792 442 1799
rect 332 1742 337 1791
rect 410 1768 417 1792
rect 355 1762 473 1768
rect 219 1738 228 1742
rect 219 1708 224 1738
rect 320 1738 337 1742
rect 248 1730 270 1734
rect 165 1688 187 1689
rect 166 1682 187 1688
rect 166 1661 172 1682
rect 251 1681 256 1730
rect 332 1689 337 1738
rect 311 1682 337 1689
rect 331 1673 337 1682
rect 80 1624 116 1632
rect 166 1563 172 1653
rect 250 1648 273 1655
rect 250 1623 257 1648
rect 225 1616 257 1623
rect 331 1622 337 1665
rect 250 1591 257 1616
rect 311 1615 337 1622
rect 192 1586 257 1591
rect 166 1556 187 1563
rect 166 1535 172 1556
rect 250 1555 257 1586
rect 331 1563 337 1615
rect 311 1556 357 1563
rect 410 1557 417 1762
rect 331 1547 337 1556
rect 166 1489 172 1527
rect 250 1522 273 1529
rect 250 1497 257 1522
rect 225 1490 257 1497
rect 331 1496 337 1539
rect 430 1529 436 1591
rect 495 1563 501 1829
rect 579 1824 602 1831
rect 579 1799 586 1824
rect 554 1792 586 1799
rect 660 1798 666 1841
rect 684 1820 688 1968
rect 579 1780 586 1792
rect 640 1791 666 1798
rect 678 1815 688 1820
rect 699 2600 725 2606
rect 779 2606 784 2638
rect 811 2628 816 2638
rect 811 2623 870 2628
rect 699 2557 705 2600
rect 779 2599 811 2606
rect 779 2574 786 2599
rect 763 2567 786 2574
rect 792 2563 798 2580
rect 864 2569 870 2623
rect 792 2559 806 2563
rect 699 2540 705 2549
rect 699 2533 725 2540
rect 699 2341 705 2533
rect 802 2451 806 2559
rect 864 2540 870 2561
rect 849 2533 870 2540
rect 864 2505 870 2533
rect 864 2499 892 2505
rect 900 2499 948 2505
rect 864 2484 871 2499
rect 802 2447 835 2451
rect 829 2374 835 2447
rect 1012 2471 1017 2675
rect 1031 2507 1036 2706
rect 1047 2538 1052 2721
rect 1063 2582 1068 3031
rect 1088 2974 1093 2988
rect 1254 2974 1259 3070
rect 1339 3005 1343 3639
rect 1290 3000 1343 3005
rect 1752 3441 1758 3832
rect 1934 3599 1962 3605
rect 1970 3599 2153 3605
rect 1934 3584 1941 3599
rect 2000 3521 2007 3546
rect 1968 3514 2095 3521
rect 1968 3498 1975 3514
rect 1934 3441 1941 3460
rect 1752 3435 1826 3441
rect 1834 3440 1941 3441
rect 2001 3440 2008 3460
rect 1834 3435 1950 3440
rect 1088 2967 1109 2974
rect 1233 2968 1259 2974
rect 1233 2967 1267 2968
rect 1088 2946 1094 2967
rect 1253 2962 1267 2967
rect 1752 2962 1758 3435
rect 1810 3415 1817 3435
rect 1877 3434 1950 3435
rect 1958 3434 2065 3440
rect 2073 3434 2123 3440
rect 1877 3415 1884 3434
rect 1934 3414 1941 3434
rect 2001 3414 2008 3434
rect 1844 3361 1851 3377
rect 2049 3414 2056 3434
rect 2116 3414 2123 3434
rect 1844 3354 1883 3361
rect 1876 3350 1883 3354
rect 1908 3350 1915 3356
rect 1968 3360 1975 3376
rect 2083 3360 2090 3376
rect 1968 3353 2053 3360
rect 2083 3353 2134 3360
rect 1876 3344 1980 3350
rect 1876 3329 1883 3344
rect 2000 3328 2007 3353
rect 2115 3328 2122 3353
rect 1810 3276 1817 3291
rect 1934 3276 1941 3290
rect 1810 3270 1838 3276
rect 1846 3275 1941 3276
rect 2049 3275 2056 3290
rect 2148 3275 2153 3599
rect 1846 3270 1962 3275
rect 1901 3127 1907 3270
rect 1934 3269 1962 3270
rect 1970 3269 2077 3275
rect 2085 3269 2153 3275
rect 2148 3128 2153 3269
rect 1934 3127 1962 3128
rect 1810 3121 1838 3127
rect 1846 3122 1962 3127
rect 1970 3122 2077 3128
rect 2085 3122 2153 3128
rect 1846 3121 1941 3122
rect 1810 3106 1817 3121
rect 1934 3107 1941 3121
rect 2049 3107 2056 3122
rect 1876 3053 1883 3068
rect 1876 3047 1980 3053
rect 1876 3043 1883 3047
rect 1844 3036 1883 3043
rect 1908 3041 1915 3047
rect 2000 3044 2007 3069
rect 2115 3044 2122 3069
rect 1968 3037 2053 3044
rect 2083 3037 2138 3044
rect 1844 3020 1851 3036
rect 1968 3021 1975 3037
rect 2083 3021 2090 3037
rect 1810 2962 1817 2982
rect 1877 2963 1884 2982
rect 1934 2963 1941 2983
rect 2001 2963 2008 2983
rect 2049 2963 2056 2983
rect 2116 2963 2123 2983
rect 1877 2962 1950 2963
rect 1253 2958 1259 2962
rect 1262 2956 1826 2962
rect 1834 2957 1950 2962
rect 1958 2957 2065 2963
rect 2073 2957 2123 2963
rect 1834 2956 1941 2957
rect 1088 2884 1094 2938
rect 1172 2933 1195 2940
rect 1172 2908 1179 2933
rect 1147 2901 1179 2908
rect 1253 2907 1259 2950
rect 1088 2879 1147 2884
rect 1088 2793 1094 2879
rect 1142 2869 1147 2879
rect 1174 2869 1179 2901
rect 1233 2901 1259 2907
rect 1934 2937 1941 2956
rect 2001 2937 2008 2957
rect 1233 2900 1260 2901
rect 1255 2869 1260 2900
rect 1968 2883 1975 2899
rect 1968 2876 2095 2883
rect 1142 2865 1151 2869
rect 1142 2835 1147 2865
rect 1243 2865 1260 2869
rect 1171 2857 1193 2861
rect 1174 2830 1179 2857
rect 1174 2825 1225 2830
rect 1089 2758 1094 2793
rect 1142 2788 1147 2803
rect 1174 2788 1179 2825
rect 1255 2788 1260 2865
rect 2000 2851 2007 2876
rect 1934 2798 1941 2813
rect 2148 2798 2153 3122
rect 1142 2784 1151 2788
rect 1142 2758 1147 2784
rect 1243 2784 1260 2788
rect 1171 2776 1193 2780
rect 1089 2754 1147 2758
rect 1089 2725 1094 2754
rect 1089 2718 1110 2725
rect 1174 2718 1179 2776
rect 1255 2768 1260 2784
rect 1464 2792 1962 2798
rect 1970 2792 2153 2798
rect 1089 2697 1095 2718
rect 1182 2751 1384 2757
rect 1182 2691 1187 2751
rect 1255 2741 1303 2745
rect 1255 2725 1260 2741
rect 1234 2718 1260 2725
rect 1254 2709 1260 2718
rect 1089 2611 1095 2689
rect 1173 2684 1196 2691
rect 1173 2659 1180 2684
rect 1148 2652 1180 2659
rect 1254 2658 1260 2701
rect 1234 2651 1260 2658
rect 1174 2615 1179 2633
rect 1142 2611 1147 2613
rect 1171 2611 1193 2615
rect 1089 2607 1147 2611
rect 1142 2603 1151 2607
rect 1255 2607 1260 2651
rect 1243 2603 1260 2607
rect 1142 2601 1147 2603
rect 1174 2582 1179 2603
rect 1255 2596 1260 2603
rect 1298 2738 1303 2741
rect 1379 2738 1384 2751
rect 1298 2734 1315 2738
rect 1298 2675 1303 2734
rect 1407 2734 1416 2738
rect 1365 2726 1387 2730
rect 1298 2668 1324 2675
rect 1379 2668 1384 2726
rect 1411 2708 1416 2734
rect 1464 2708 1469 2792
rect 1411 2704 1469 2708
rect 1464 2675 1469 2704
rect 1448 2668 1469 2675
rect 1298 2659 1304 2668
rect 1298 2608 1304 2651
rect 1463 2647 1469 2668
rect 1362 2634 1385 2641
rect 1378 2609 1385 2634
rect 1298 2601 1324 2608
rect 1378 2602 1410 2609
rect 1063 2576 1179 2582
rect 1148 2571 1153 2576
rect 1298 2557 1303 2601
rect 1378 2597 1385 2602
rect 1463 2601 1469 2639
rect 1379 2565 1384 2583
rect 1365 2561 1387 2565
rect 1411 2561 1416 2563
rect 1464 2561 1469 2601
rect 1298 2553 1315 2557
rect 1411 2557 1469 2561
rect 1407 2553 1416 2557
rect 1298 2546 1303 2553
rect 1379 2538 1384 2553
rect 1411 2551 1416 2553
rect 1047 2534 1384 2538
rect 1305 2526 1311 2534
rect 1031 2502 1366 2507
rect 1012 2467 1343 2471
rect 930 2421 937 2446
rect 898 2414 1025 2421
rect 898 2398 905 2414
rect 864 2341 871 2360
rect 699 2335 756 2341
rect 764 2340 871 2341
rect 931 2340 938 2360
rect 1167 2340 1217 2341
rect 764 2335 880 2340
rect 699 1956 705 2335
rect 740 2315 747 2335
rect 807 2334 880 2335
rect 888 2334 995 2340
rect 1003 2334 1110 2340
rect 1118 2336 1217 2340
rect 1118 2334 1168 2336
rect 807 2315 814 2334
rect 864 2314 871 2334
rect 931 2314 938 2334
rect 774 2261 781 2277
rect 979 2314 986 2334
rect 1046 2314 1053 2334
rect 1094 2314 1101 2334
rect 1161 2314 1168 2334
rect 1199 2324 1203 2336
rect 774 2254 813 2261
rect 806 2250 813 2254
rect 838 2250 845 2256
rect 898 2260 905 2276
rect 1013 2260 1020 2276
rect 1128 2260 1135 2276
rect 1207 2260 1211 2274
rect 1313 2260 1318 2410
rect 898 2253 983 2260
rect 1013 2253 1066 2260
rect 806 2244 910 2250
rect 806 2229 813 2244
rect 930 2228 937 2253
rect 1045 2252 1066 2253
rect 1128 2255 1199 2260
rect 1207 2255 1331 2260
rect 1128 2253 1167 2255
rect 1045 2228 1052 2252
rect 1160 2228 1167 2253
rect 1207 2252 1211 2255
rect 1199 2228 1203 2232
rect 740 2176 747 2191
rect 1184 2223 1213 2228
rect 864 2176 871 2190
rect 740 2170 768 2176
rect 776 2175 871 2176
rect 979 2175 986 2190
rect 1094 2175 1101 2190
rect 1184 2175 1189 2223
rect 776 2170 892 2175
rect 864 2169 892 2170
rect 900 2169 1007 2175
rect 1015 2169 1122 2175
rect 1130 2169 1189 2175
rect 1072 2122 1077 2169
rect 864 2121 892 2122
rect 740 2115 768 2121
rect 776 2116 892 2121
rect 900 2116 1007 2122
rect 1015 2116 1077 2122
rect 1094 2154 1101 2169
rect 1184 2121 1189 2169
rect 1184 2116 1213 2121
rect 776 2115 871 2116
rect 740 2100 747 2115
rect 864 2101 871 2115
rect 979 2101 986 2116
rect 1160 2091 1167 2116
rect 1199 2112 1203 2116
rect 1128 2089 1167 2091
rect 1207 2089 1211 2092
rect 1313 2089 1317 2175
rect 1128 2084 1199 2089
rect 1207 2084 1317 2089
rect 1128 2068 1135 2084
rect 1207 2070 1211 2084
rect 806 2047 813 2062
rect 806 2041 910 2047
rect 806 2037 813 2041
rect 774 2030 813 2037
rect 838 2035 845 2041
rect 930 2038 937 2063
rect 1045 2039 1052 2063
rect 1045 2038 1066 2039
rect 898 2031 983 2038
rect 1013 2031 1066 2038
rect 774 2014 781 2030
rect 898 2015 905 2031
rect 1013 2015 1020 2031
rect 740 1956 747 1976
rect 807 1957 814 1976
rect 864 1957 871 1977
rect 931 1957 938 1977
rect 1094 2010 1101 2030
rect 1161 2010 1168 2030
rect 1094 2004 1110 2010
rect 1118 2009 1168 2010
rect 1199 2009 1203 2020
rect 1118 2004 1217 2009
rect 1094 1994 1101 2004
rect 1192 2003 1217 2004
rect 1167 1994 1217 1995
rect 979 1957 986 1977
rect 1046 1957 1053 1977
rect 1068 1989 1110 1994
rect 1068 1957 1073 1989
rect 807 1956 880 1957
rect 699 1950 756 1956
rect 764 1951 880 1956
rect 888 1951 995 1957
rect 1003 1951 1073 1957
rect 1094 1988 1110 1989
rect 1118 1990 1217 1994
rect 1118 1988 1168 1990
rect 1094 1968 1101 1988
rect 1161 1968 1168 1988
rect 764 1950 871 1951
rect 481 1556 502 1563
rect 395 1522 436 1529
rect 496 1535 502 1556
rect 411 1497 418 1522
rect 250 1469 257 1490
rect 311 1489 357 1496
rect 411 1490 443 1497
rect 496 1494 502 1527
rect 678 1512 682 1815
rect 699 1758 705 1950
rect 864 1931 871 1950
rect 931 1931 938 1951
rect 829 1844 835 1917
rect 1199 1978 1203 1990
rect 1128 1914 1135 1930
rect 1228 1941 1233 2084
rect 1326 1978 1331 2255
rect 1241 1974 1331 1978
rect 1339 2172 1343 2467
rect 1361 2383 1366 2502
rect 1464 2409 1469 2557
rect 2148 2479 2153 2792
rect 1934 2473 1962 2479
rect 1970 2473 2153 2479
rect 1934 2458 1941 2473
rect 1464 2405 1479 2409
rect 1474 2383 1479 2405
rect 2000 2395 2007 2420
rect 1361 2379 1378 2383
rect 1470 2379 1479 2383
rect 1361 2320 1366 2379
rect 1428 2371 1450 2375
rect 1361 2313 1387 2320
rect 1442 2313 1447 2371
rect 1474 2353 1479 2379
rect 1968 2388 2095 2395
rect 1968 2372 1975 2388
rect 1474 2349 1532 2353
rect 1527 2320 1532 2349
rect 1511 2313 1532 2320
rect 1934 2315 1941 2334
rect 1361 2304 1367 2313
rect 1361 2253 1367 2296
rect 1526 2292 1532 2313
rect 1425 2279 1448 2286
rect 1441 2254 1448 2279
rect 1361 2246 1387 2253
rect 1441 2247 1473 2254
rect 1361 2202 1366 2246
rect 1441 2243 1448 2247
rect 1526 2246 1532 2284
rect 1442 2210 1447 2228
rect 1428 2206 1450 2210
rect 1474 2206 1479 2208
rect 1527 2206 1532 2246
rect 1706 2309 1826 2315
rect 1834 2314 1941 2315
rect 2001 2314 2008 2334
rect 1834 2309 1950 2314
rect 1706 2213 1711 2309
rect 1810 2289 1817 2309
rect 1877 2308 1950 2309
rect 1958 2308 2065 2314
rect 2073 2308 2123 2314
rect 1877 2289 1884 2308
rect 1934 2288 1941 2308
rect 2001 2288 2008 2308
rect 1844 2235 1851 2251
rect 2049 2288 2056 2308
rect 2116 2288 2123 2308
rect 1844 2228 1883 2235
rect 1474 2202 1532 2206
rect 1361 2198 1378 2202
rect 1470 2198 1479 2202
rect 1339 2168 1352 2172
rect 1241 1973 1246 1974
rect 1228 1936 1268 1941
rect 1207 1914 1211 1928
rect 1128 1909 1199 1914
rect 1207 1909 1283 1914
rect 1128 1907 1167 1909
rect 898 1877 905 1893
rect 1160 1882 1167 1907
rect 1207 1906 1211 1909
rect 1199 1882 1203 1886
rect 898 1870 1025 1877
rect 930 1845 937 1870
rect 802 1840 835 1844
rect 699 1751 725 1758
rect 699 1742 705 1751
rect 699 1691 705 1734
rect 802 1732 806 1840
rect 1184 1877 1213 1882
rect 1094 1829 1101 1844
rect 1184 1829 1189 1877
rect 1094 1823 1122 1829
rect 1130 1823 1189 1829
rect 864 1792 871 1807
rect 1094 1792 1101 1823
rect 864 1786 892 1792
rect 900 1787 1119 1792
rect 900 1786 1077 1787
rect 1091 1786 1119 1787
rect 1127 1786 1186 1792
rect 864 1758 870 1786
rect 849 1751 870 1758
rect 792 1728 806 1732
rect 864 1730 870 1751
rect 1091 1771 1098 1786
rect 1181 1738 1186 1786
rect 1181 1733 1211 1738
rect 763 1717 786 1724
rect 779 1692 786 1717
rect 792 1711 798 1728
rect 699 1685 725 1691
rect 698 1684 725 1685
rect 779 1685 811 1692
rect 698 1653 703 1684
rect 779 1653 784 1685
rect 864 1668 870 1722
rect 1157 1708 1164 1733
rect 1196 1729 1200 1733
rect 1339 1717 1343 2168
rect 1361 2166 1366 2198
rect 1474 2196 1479 2198
rect 1361 2163 1370 2166
rect 1365 2148 1370 2163
rect 1527 2157 1532 2202
rect 1593 2209 1602 2213
rect 1694 2209 1711 2213
rect 1593 2183 1598 2209
rect 1622 2201 1644 2205
rect 1540 2179 1598 2183
rect 1540 2157 1545 2179
rect 1527 2151 1545 2157
rect 1365 2144 1382 2148
rect 1474 2144 1483 2148
rect 1365 2085 1370 2144
rect 1432 2136 1454 2140
rect 1365 2078 1391 2085
rect 1446 2078 1451 2136
rect 1478 2118 1483 2144
rect 1531 2118 1536 2151
rect 1478 2114 1536 2118
rect 1531 2085 1536 2114
rect 1515 2078 1536 2085
rect 1365 2069 1371 2078
rect 1365 2018 1371 2061
rect 1530 2057 1536 2078
rect 1429 2044 1452 2051
rect 1445 2019 1452 2044
rect 1365 2011 1391 2018
rect 1445 2012 1477 2019
rect 1365 1967 1370 2011
rect 1445 2007 1452 2012
rect 1530 2011 1536 2049
rect 1540 2150 1545 2151
rect 1540 2143 1561 2150
rect 1625 2143 1630 2201
rect 1540 2122 1546 2143
rect 1633 2165 1640 2170
rect 1633 2116 1637 2165
rect 1706 2150 1711 2209
rect 1876 2224 1883 2228
rect 1908 2224 1915 2230
rect 1968 2234 1975 2250
rect 2083 2234 2090 2250
rect 1968 2227 2053 2234
rect 2083 2227 2136 2234
rect 1876 2218 1980 2224
rect 1876 2203 1883 2218
rect 1685 2143 1711 2150
rect 2000 2202 2007 2227
rect 2115 2202 2122 2227
rect 1810 2150 1817 2165
rect 1934 2150 1941 2164
rect 1810 2144 1838 2150
rect 1846 2149 1941 2150
rect 2049 2149 2056 2164
rect 2148 2149 2153 2473
rect 1846 2144 1962 2149
rect 1934 2143 1962 2144
rect 1970 2143 2077 2149
rect 2085 2143 2153 2149
rect 1705 2134 1711 2143
rect 1540 2076 1546 2114
rect 1624 2109 1647 2116
rect 1624 2084 1631 2109
rect 1599 2077 1631 2084
rect 1705 2083 1711 2126
rect 1540 2036 1545 2076
rect 1624 2072 1631 2077
rect 1685 2076 1711 2083
rect 1625 2040 1630 2058
rect 1593 2036 1598 2038
rect 1622 2036 1644 2040
rect 1540 2032 1598 2036
rect 1706 2032 1711 2076
rect 1593 2028 1602 2032
rect 1694 2028 1711 2032
rect 1593 2026 1598 2028
rect 1446 1975 1451 1993
rect 1432 1971 1454 1975
rect 1478 1971 1483 1973
rect 1531 1971 1536 2011
rect 1478 1967 1536 1971
rect 1365 1963 1382 1967
rect 1474 1963 1483 1967
rect 1365 1735 1370 1963
rect 1478 1961 1483 1963
rect 1531 1737 1536 1967
rect 1706 1836 1711 2028
rect 2148 2002 2153 2143
rect 1934 2001 1962 2002
rect 1810 1995 1838 2001
rect 1846 1996 1962 2001
rect 1970 1996 2077 2002
rect 2085 1996 2153 2002
rect 1846 1995 1941 1996
rect 1810 1980 1817 1995
rect 1934 1981 1941 1995
rect 2049 1981 2056 1996
rect 1876 1927 1883 1942
rect 1876 1921 1980 1927
rect 1876 1917 1883 1921
rect 1844 1910 1883 1917
rect 1908 1915 1915 1921
rect 2000 1918 2007 1943
rect 2115 1918 2122 1943
rect 1968 1911 2053 1918
rect 2083 1911 2138 1918
rect 1844 1894 1851 1910
rect 1968 1895 1975 1911
rect 2083 1895 2090 1911
rect 1810 1836 1817 1856
rect 1877 1837 1884 1856
rect 1934 1837 1941 1857
rect 2001 1837 2008 1857
rect 2049 1837 2056 1857
rect 2116 1837 2123 1857
rect 1877 1836 1950 1837
rect 1706 1830 1826 1836
rect 1834 1831 1950 1836
rect 1958 1831 2065 1837
rect 2073 1831 2123 1837
rect 1834 1830 1941 1831
rect 1934 1811 1941 1830
rect 2001 1811 2008 1831
rect 1968 1757 1975 1773
rect 1968 1750 2095 1757
rect 1365 1731 1463 1735
rect 1531 1733 1576 1737
rect 1125 1706 1164 1708
rect 1204 1706 1208 1709
rect 1125 1701 1196 1706
rect 1204 1701 1395 1706
rect 1125 1685 1132 1701
rect 1204 1687 1208 1701
rect 811 1663 870 1668
rect 811 1653 816 1663
rect 698 1649 715 1653
rect 698 1585 703 1649
rect 807 1649 816 1653
rect 765 1641 787 1645
rect 779 1601 784 1641
rect 811 1624 816 1649
rect 1091 1627 1098 1647
rect 1158 1627 1165 1647
rect 811 1619 1075 1624
rect 1091 1621 1107 1627
rect 1115 1625 1165 1627
rect 1196 1625 1200 1637
rect 1458 1625 1463 1731
rect 1115 1621 1463 1625
rect 1164 1620 1463 1621
rect 779 1595 1061 1601
rect 698 1580 1033 1585
rect 678 1507 999 1512
rect 678 1494 682 1507
rect 250 1463 303 1469
rect 331 1442 337 1489
rect 411 1466 418 1490
rect 496 1489 682 1494
rect 0 1436 666 1442
rect 0 1386 6 1436
rect 165 1411 501 1417
rect 0 1379 26 1386
rect 0 1370 6 1379
rect 0 1319 6 1362
rect 80 1352 87 1388
rect 165 1386 171 1411
rect 495 1386 501 1411
rect 660 1386 666 1436
rect 150 1379 186 1386
rect 310 1379 356 1386
rect 480 1379 516 1386
rect 640 1379 666 1386
rect 64 1345 87 1352
rect 80 1320 87 1345
rect 165 1358 171 1379
rect 330 1370 336 1379
rect 0 1312 26 1319
rect 80 1313 112 1320
rect 0 963 6 1312
rect 80 1153 87 1313
rect 165 1278 171 1350
rect 249 1345 272 1352
rect 249 1320 256 1345
rect 224 1313 256 1320
rect 330 1319 336 1362
rect 495 1358 501 1379
rect 394 1345 417 1352
rect 410 1320 417 1345
rect 660 1370 666 1379
rect 165 1273 224 1278
rect 165 1210 171 1273
rect 219 1263 224 1273
rect 251 1263 256 1313
rect 310 1312 356 1319
rect 410 1313 442 1320
rect 332 1263 337 1312
rect 410 1289 417 1313
rect 355 1283 473 1289
rect 219 1259 228 1263
rect 219 1229 224 1259
rect 320 1259 337 1263
rect 248 1251 270 1255
rect 165 1209 187 1210
rect 166 1203 187 1209
rect 166 1182 172 1203
rect 251 1202 256 1251
rect 332 1210 337 1259
rect 311 1203 337 1210
rect 331 1194 337 1203
rect 80 1145 116 1153
rect 166 1084 172 1174
rect 250 1169 273 1176
rect 250 1144 257 1169
rect 225 1137 257 1144
rect 331 1143 337 1186
rect 250 1112 257 1137
rect 311 1136 337 1143
rect 192 1107 257 1112
rect 166 1077 187 1084
rect 166 1056 172 1077
rect 250 1076 257 1107
rect 331 1084 337 1136
rect 311 1077 357 1084
rect 410 1078 417 1283
rect 331 1068 337 1077
rect 166 1010 172 1048
rect 250 1043 273 1050
rect 250 1018 257 1043
rect 225 1011 257 1018
rect 331 1017 337 1060
rect 430 1050 436 1112
rect 495 1084 501 1350
rect 579 1345 602 1352
rect 579 1320 586 1345
rect 554 1313 586 1320
rect 660 1319 666 1362
rect 579 1301 586 1313
rect 640 1312 666 1319
rect 481 1077 502 1084
rect 395 1043 436 1050
rect 496 1056 502 1077
rect 411 1018 418 1043
rect 250 990 257 1011
rect 311 1010 357 1017
rect 411 1011 443 1018
rect 496 1015 502 1048
rect 678 1015 682 1489
rect 250 984 303 990
rect 331 963 337 1010
rect 411 987 418 1011
rect 496 1010 682 1015
rect 0 957 666 963
rect 0 907 6 957
rect 165 932 501 938
rect 0 900 26 907
rect 0 891 6 900
rect 0 840 6 883
rect 80 873 87 909
rect 165 907 171 932
rect 495 907 501 932
rect 660 907 666 957
rect 150 900 186 907
rect 310 900 356 907
rect 480 900 516 907
rect 640 900 666 907
rect 64 866 87 873
rect 80 841 87 866
rect 165 879 171 900
rect 330 891 336 900
rect 0 833 26 840
rect 80 834 112 841
rect 0 484 6 833
rect 80 674 87 834
rect 165 799 171 871
rect 249 866 272 873
rect 249 841 256 866
rect 224 834 256 841
rect 330 840 336 883
rect 495 879 501 900
rect 394 866 417 873
rect 410 841 417 866
rect 660 891 666 900
rect 165 794 224 799
rect 165 731 171 794
rect 219 784 224 794
rect 251 784 256 834
rect 310 833 356 840
rect 410 834 442 841
rect 332 784 337 833
rect 410 810 417 834
rect 355 804 473 810
rect 219 780 228 784
rect 219 750 224 780
rect 320 780 337 784
rect 248 772 270 776
rect 165 730 187 731
rect 166 724 187 730
rect 166 703 172 724
rect 251 723 256 772
rect 332 731 337 780
rect 311 724 337 731
rect 331 715 337 724
rect 80 666 116 674
rect 166 605 172 695
rect 250 690 273 697
rect 250 665 257 690
rect 225 658 257 665
rect 331 664 337 707
rect 250 633 257 658
rect 311 657 337 664
rect 192 628 257 633
rect 166 598 187 605
rect 166 577 172 598
rect 250 597 257 628
rect 331 605 337 657
rect 311 598 357 605
rect 410 599 417 804
rect 331 589 337 598
rect 166 531 172 569
rect 250 564 273 571
rect 250 539 257 564
rect 225 532 257 539
rect 331 538 337 581
rect 430 571 436 633
rect 495 605 501 871
rect 579 866 602 873
rect 579 841 586 866
rect 554 834 586 841
rect 660 840 666 883
rect 579 822 586 834
rect 640 833 666 840
rect 481 598 502 605
rect 395 564 436 571
rect 496 577 502 598
rect 411 539 418 564
rect 250 511 257 532
rect 311 531 357 538
rect 411 532 443 539
rect 496 536 502 569
rect 678 536 682 1010
rect 994 958 999 1507
rect 1028 1419 1033 1580
rect 1056 1443 1061 1595
rect 1070 1591 1075 1619
rect 1458 1612 1463 1620
rect 1571 1612 1576 1733
rect 2000 1725 2007 1750
rect 1934 1672 1941 1687
rect 2148 1672 2153 1996
rect 1934 1671 1962 1672
rect 1458 1608 1475 1612
rect 1567 1608 1576 1612
rect 1070 1586 1115 1591
rect 1087 1585 1115 1586
rect 1123 1585 1182 1591
rect 1087 1570 1094 1585
rect 1177 1537 1182 1585
rect 1458 1549 1463 1608
rect 1525 1600 1547 1604
rect 1458 1542 1484 1549
rect 1539 1542 1544 1600
rect 1571 1582 1576 1608
rect 1624 1666 1962 1671
rect 1970 1666 2153 1672
rect 2177 3275 2183 3832
rect 2299 3823 2306 3848
rect 2233 3770 2240 3785
rect 2535 3770 2563 3771
rect 2202 3764 2261 3770
rect 2269 3765 2563 3770
rect 2571 3765 2679 3771
rect 2269 3764 2542 3765
rect 2202 3440 2208 3764
rect 2233 3749 2240 3764
rect 2535 3750 2542 3764
rect 2299 3686 2306 3711
rect 2330 3686 2336 3742
rect 2601 3687 2608 3712
rect 2267 3679 2541 3686
rect 2569 3680 2632 3687
rect 2267 3663 2274 3679
rect 2233 3605 2240 3625
rect 2300 3606 2307 3625
rect 2330 3624 2336 3679
rect 2569 3664 2576 3680
rect 2535 3606 2542 3626
rect 2602 3606 2609 3626
rect 2300 3605 2425 3606
rect 2233 3599 2249 3605
rect 2257 3601 2425 3605
rect 2257 3599 2307 3601
rect 2233 3579 2240 3599
rect 2300 3579 2307 3599
rect 2356 3589 2360 3601
rect 2409 3600 2425 3601
rect 2433 3600 2551 3606
rect 2559 3600 2661 3606
rect 2267 3525 2274 3541
rect 2409 3580 2416 3600
rect 2476 3580 2483 3600
rect 2535 3580 2542 3600
rect 2602 3580 2609 3600
rect 2364 3525 2368 3539
rect 2443 3526 2450 3542
rect 2569 3526 2576 3542
rect 2629 3526 2635 3572
rect 2267 3520 2356 3525
rect 2364 3520 2417 3525
rect 2267 3518 2306 3520
rect 2299 3493 2306 3518
rect 2364 3517 2368 3520
rect 2443 3519 2543 3526
rect 2569 3519 2635 3526
rect 2356 3493 2360 3497
rect 2475 3494 2482 3519
rect 2341 3488 2390 3493
rect 2233 3440 2240 3455
rect 2341 3440 2346 3488
rect 2507 3461 2512 3519
rect 2601 3494 2608 3519
rect 2409 3441 2416 3456
rect 2535 3441 2542 3456
rect 2409 3440 2437 3441
rect 2202 3434 2261 3440
rect 2269 3435 2437 3440
rect 2445 3435 2563 3441
rect 2571 3435 2609 3441
rect 2269 3434 2410 3435
rect 2233 3419 2240 3434
rect 2299 3356 2306 3381
rect 2466 3356 2474 3385
rect 2231 3349 2474 3356
rect 2267 3333 2274 3349
rect 2233 3275 2240 3295
rect 2300 3275 2307 3295
rect 2656 3275 2661 3600
rect 2177 3269 2249 3275
rect 2257 3269 2661 3275
rect 2177 2615 2183 3269
rect 2233 3249 2240 3269
rect 2300 3249 2307 3269
rect 2267 3195 2274 3211
rect 2267 3188 2318 3195
rect 2299 3163 2306 3188
rect 2233 3110 2240 3125
rect 2674 3111 2679 3765
rect 2535 3110 2563 3111
rect 2202 3104 2261 3110
rect 2269 3105 2563 3110
rect 2571 3105 2679 3111
rect 2269 3104 2542 3105
rect 2202 2780 2208 3104
rect 2233 3089 2240 3104
rect 2535 3090 2542 3104
rect 2299 3026 2306 3051
rect 2330 3026 2336 3082
rect 2601 3027 2608 3052
rect 2267 3019 2541 3026
rect 2569 3020 2632 3027
rect 2267 3003 2274 3019
rect 2233 2945 2240 2965
rect 2300 2946 2307 2965
rect 2330 2964 2336 3019
rect 2569 3004 2576 3020
rect 2535 2946 2542 2966
rect 2602 2946 2609 2966
rect 2300 2945 2425 2946
rect 2233 2939 2249 2945
rect 2257 2941 2425 2945
rect 2257 2939 2307 2941
rect 2233 2919 2240 2939
rect 2300 2919 2307 2939
rect 2356 2929 2360 2941
rect 2409 2940 2425 2941
rect 2433 2940 2551 2946
rect 2559 2940 2661 2946
rect 2267 2865 2274 2881
rect 2409 2920 2416 2940
rect 2476 2920 2483 2940
rect 2535 2920 2542 2940
rect 2602 2920 2609 2940
rect 2364 2865 2368 2879
rect 2443 2866 2450 2882
rect 2569 2866 2576 2882
rect 2629 2866 2635 2912
rect 2267 2860 2356 2865
rect 2364 2860 2417 2865
rect 2267 2858 2306 2860
rect 2299 2833 2306 2858
rect 2364 2857 2368 2860
rect 2443 2859 2543 2866
rect 2569 2859 2635 2866
rect 2356 2833 2360 2837
rect 2475 2834 2482 2859
rect 2341 2828 2390 2833
rect 2233 2780 2240 2795
rect 2341 2780 2346 2828
rect 2507 2801 2512 2859
rect 2601 2834 2608 2859
rect 2409 2781 2416 2796
rect 2535 2781 2542 2796
rect 2409 2780 2437 2781
rect 2202 2774 2261 2780
rect 2269 2775 2437 2780
rect 2445 2775 2563 2781
rect 2571 2775 2609 2781
rect 2269 2774 2410 2775
rect 2233 2759 2240 2774
rect 2299 2696 2306 2721
rect 2466 2696 2474 2725
rect 2231 2689 2474 2696
rect 2267 2673 2274 2689
rect 2233 2615 2240 2635
rect 2300 2615 2307 2635
rect 2656 2615 2661 2940
rect 2177 2609 2249 2615
rect 2257 2609 2661 2615
rect 2177 1955 2183 2609
rect 2233 2589 2240 2609
rect 2300 2589 2307 2609
rect 2267 2535 2274 2551
rect 2267 2528 2318 2535
rect 2299 2503 2306 2528
rect 2233 2450 2240 2465
rect 2674 2451 2679 3105
rect 2535 2450 2563 2451
rect 2202 2444 2261 2450
rect 2269 2445 2563 2450
rect 2571 2445 2679 2451
rect 2269 2444 2542 2445
rect 2202 2120 2208 2444
rect 2233 2429 2240 2444
rect 2535 2430 2542 2444
rect 2299 2366 2306 2391
rect 2330 2366 2336 2422
rect 2601 2367 2608 2392
rect 2267 2359 2541 2366
rect 2569 2360 2632 2367
rect 2267 2343 2274 2359
rect 2233 2285 2240 2305
rect 2300 2286 2307 2305
rect 2330 2304 2336 2359
rect 2569 2344 2576 2360
rect 2535 2286 2542 2306
rect 2602 2286 2609 2306
rect 2300 2285 2425 2286
rect 2233 2279 2249 2285
rect 2257 2281 2425 2285
rect 2257 2279 2307 2281
rect 2233 2259 2240 2279
rect 2300 2259 2307 2279
rect 2356 2269 2360 2281
rect 2409 2280 2425 2281
rect 2433 2280 2551 2286
rect 2559 2280 2661 2286
rect 2267 2205 2274 2221
rect 2409 2260 2416 2280
rect 2476 2260 2483 2280
rect 2535 2260 2542 2280
rect 2602 2260 2609 2280
rect 2364 2205 2368 2219
rect 2443 2206 2450 2222
rect 2569 2206 2576 2222
rect 2629 2206 2635 2252
rect 2267 2200 2356 2205
rect 2364 2200 2417 2205
rect 2267 2198 2306 2200
rect 2299 2173 2306 2198
rect 2364 2197 2368 2200
rect 2443 2199 2543 2206
rect 2569 2199 2635 2206
rect 2356 2173 2360 2177
rect 2475 2174 2482 2199
rect 2341 2168 2390 2173
rect 2233 2120 2240 2135
rect 2341 2120 2346 2168
rect 2507 2141 2512 2199
rect 2601 2174 2608 2199
rect 2409 2121 2416 2136
rect 2535 2121 2542 2136
rect 2409 2120 2437 2121
rect 2202 2114 2261 2120
rect 2269 2115 2437 2120
rect 2445 2115 2563 2121
rect 2571 2115 2609 2121
rect 2269 2114 2410 2115
rect 2233 2099 2240 2114
rect 2299 2036 2306 2061
rect 2466 2036 2474 2065
rect 2231 2029 2474 2036
rect 2267 2013 2274 2029
rect 2233 1955 2240 1975
rect 2300 1955 2307 1975
rect 2656 1955 2661 2280
rect 2177 1949 2249 1955
rect 2257 1949 2661 1955
rect 1624 1582 1629 1666
rect 1571 1578 1629 1582
rect 1624 1549 1629 1578
rect 1608 1542 1629 1549
rect 1177 1532 1205 1537
rect 1458 1533 1464 1542
rect 1153 1507 1160 1532
rect 1192 1528 1196 1532
rect 1121 1505 1160 1507
rect 1200 1505 1204 1508
rect 1121 1500 1192 1505
rect 1200 1500 1431 1505
rect 1121 1484 1128 1500
rect 1200 1486 1204 1500
rect 1087 1426 1094 1446
rect 1154 1426 1161 1446
rect 1087 1420 1103 1426
rect 1111 1424 1161 1426
rect 1192 1424 1196 1436
rect 1111 1420 1215 1424
rect 1087 1419 1093 1420
rect 1160 1419 1215 1420
rect 1425 1420 1431 1500
rect 1028 1413 1093 1419
rect 1458 1482 1464 1525
rect 1623 1521 1629 1542
rect 1522 1508 1545 1515
rect 1538 1483 1545 1508
rect 1458 1475 1484 1482
rect 1538 1476 1570 1483
rect 1458 1431 1463 1475
rect 1538 1472 1545 1476
rect 1623 1475 1629 1513
rect 1539 1439 1544 1457
rect 1525 1435 1547 1439
rect 1571 1435 1576 1437
rect 1624 1435 1629 1475
rect 1803 1442 1808 1449
rect 1571 1431 1629 1435
rect 1458 1427 1475 1431
rect 1567 1427 1576 1431
rect 1028 1011 1033 1413
rect 1087 1412 1093 1413
rect 1160 1412 1215 1413
rect 1087 1406 1103 1412
rect 1111 1408 1215 1412
rect 1111 1406 1161 1408
rect 1087 1386 1094 1406
rect 1154 1386 1161 1406
rect 1192 1396 1196 1408
rect 1121 1332 1128 1348
rect 1200 1332 1204 1346
rect 1442 1332 1448 1401
rect 1458 1394 1463 1427
rect 1571 1425 1576 1427
rect 1624 1419 1629 1431
rect 1690 1438 1699 1442
rect 1791 1438 1808 1442
rect 1690 1419 1695 1438
rect 1719 1430 1741 1434
rect 1624 1415 1695 1419
rect 1624 1414 1642 1415
rect 1458 1389 1467 1394
rect 1121 1327 1192 1332
rect 1200 1327 1448 1332
rect 1462 1377 1467 1389
rect 1637 1379 1642 1414
rect 1462 1373 1479 1377
rect 1571 1373 1580 1377
rect 1121 1325 1160 1327
rect 1153 1300 1160 1325
rect 1200 1324 1204 1327
rect 1462 1314 1467 1373
rect 1529 1365 1551 1369
rect 1462 1307 1488 1314
rect 1543 1307 1548 1365
rect 1575 1347 1580 1373
rect 1628 1372 1658 1379
rect 1722 1372 1727 1430
rect 1628 1347 1633 1372
rect 1575 1343 1633 1347
rect 1628 1314 1633 1343
rect 1612 1307 1633 1314
rect 1192 1300 1196 1304
rect 1177 1295 1225 1300
rect 1462 1298 1468 1307
rect 1087 1247 1094 1262
rect 1177 1247 1182 1295
rect 1087 1246 1115 1247
rect 1077 1241 1115 1246
rect 1123 1246 1182 1247
rect 1462 1247 1468 1290
rect 1627 1286 1633 1307
rect 1526 1273 1549 1280
rect 1542 1248 1549 1273
rect 1123 1241 1192 1246
rect 1077 1218 1082 1241
rect 1462 1240 1488 1247
rect 1542 1241 1574 1248
rect 1077 1213 1115 1218
rect 1087 1212 1115 1213
rect 1123 1213 1192 1218
rect 1123 1212 1182 1213
rect 1087 1197 1094 1212
rect 1177 1164 1182 1212
rect 1462 1196 1467 1240
rect 1542 1236 1549 1241
rect 1627 1240 1633 1278
rect 1637 1351 1643 1372
rect 1730 1400 1750 1404
rect 1730 1345 1735 1400
rect 1803 1379 1808 1438
rect 1782 1372 1808 1379
rect 1802 1363 1808 1372
rect 1637 1265 1643 1343
rect 1721 1338 1744 1345
rect 1721 1313 1728 1338
rect 1696 1306 1728 1313
rect 1802 1312 1808 1355
rect 1721 1301 1728 1306
rect 1782 1305 1808 1312
rect 1722 1269 1727 1287
rect 1690 1265 1695 1267
rect 1719 1265 1741 1269
rect 1637 1261 1695 1265
rect 1803 1261 1808 1305
rect 1690 1257 1699 1261
rect 1791 1257 1808 1261
rect 1690 1255 1695 1257
rect 1803 1241 1808 1257
rect 1543 1204 1548 1222
rect 1529 1200 1551 1204
rect 1575 1200 1580 1202
rect 1628 1200 1633 1240
rect 1575 1196 1633 1200
rect 1462 1192 1479 1196
rect 1571 1192 1580 1196
rect 1177 1159 1225 1164
rect 1153 1134 1160 1159
rect 1192 1155 1196 1159
rect 1121 1132 1160 1134
rect 1200 1132 1204 1135
rect 1121 1127 1192 1132
rect 1200 1127 1419 1132
rect 1121 1111 1128 1127
rect 1200 1113 1204 1127
rect 1087 1053 1094 1073
rect 1154 1053 1161 1073
rect 1087 1047 1103 1053
rect 1111 1051 1161 1053
rect 1192 1051 1196 1063
rect 1111 1047 1215 1051
rect 1087 1011 1093 1047
rect 1160 1046 1215 1047
rect 1462 1011 1467 1192
rect 1575 1190 1580 1192
rect 1028 1006 1467 1011
rect 1628 1150 1633 1196
rect 1794 1236 1808 1241
rect 1681 1180 1686 1191
rect 1794 1180 1799 1236
rect 1681 1176 1690 1180
rect 1782 1176 1799 1180
rect 1681 1150 1686 1176
rect 1710 1168 1732 1172
rect 1628 1146 1686 1150
rect 1628 1117 1633 1146
rect 1628 1110 1649 1117
rect 1713 1110 1718 1168
rect 1628 1089 1634 1110
rect 1721 1083 1725 1148
rect 1794 1117 1799 1176
rect 1773 1110 1799 1117
rect 1793 1101 1799 1110
rect 1628 1043 1634 1081
rect 1712 1076 1735 1083
rect 1712 1051 1719 1076
rect 1687 1044 1719 1051
rect 1793 1050 1799 1093
rect 1628 1003 1633 1043
rect 1712 1039 1719 1044
rect 1773 1043 1799 1050
rect 1713 1007 1718 1025
rect 1681 1003 1686 1005
rect 1710 1003 1732 1007
rect 1628 999 1686 1003
rect 1794 999 1799 1043
rect 1628 958 1633 999
rect 1681 995 1690 999
rect 1782 995 1799 999
rect 1681 993 1686 995
rect 994 953 1633 958
rect 1794 941 1799 995
rect 250 505 303 511
rect 331 484 337 531
rect 411 508 418 532
rect 496 531 682 536
rect 0 478 666 484
rect 0 428 6 478
rect 165 453 501 459
rect 0 421 26 428
rect 0 412 6 421
rect 0 361 6 404
rect 80 394 87 430
rect 165 428 171 453
rect 495 428 501 453
rect 660 428 666 478
rect 150 421 186 428
rect 310 421 356 428
rect 480 421 516 428
rect 640 421 666 428
rect 64 387 87 394
rect 80 362 87 387
rect 165 400 171 421
rect 330 412 336 421
rect 0 354 26 361
rect 80 355 112 362
rect 0 5 6 354
rect 80 195 87 355
rect 165 320 171 392
rect 249 387 272 394
rect 249 362 256 387
rect 224 355 256 362
rect 330 361 336 404
rect 495 400 501 421
rect 394 387 417 394
rect 410 362 417 387
rect 660 412 666 421
rect 165 315 224 320
rect 165 252 171 315
rect 219 305 224 315
rect 251 305 256 355
rect 310 354 356 361
rect 410 355 442 362
rect 332 305 337 354
rect 410 331 417 355
rect 355 325 473 331
rect 219 301 228 305
rect 219 271 224 301
rect 320 301 337 305
rect 248 293 270 297
rect 165 251 187 252
rect 166 245 187 251
rect 166 224 172 245
rect 251 244 256 293
rect 332 252 337 301
rect 311 245 337 252
rect 331 236 337 245
rect 80 187 116 195
rect 166 126 172 216
rect 250 211 273 218
rect 250 186 257 211
rect 225 179 257 186
rect 331 185 337 228
rect 250 154 257 179
rect 311 178 337 185
rect 192 149 257 154
rect 166 119 187 126
rect 166 98 172 119
rect 250 118 257 149
rect 331 126 337 178
rect 311 119 357 126
rect 410 120 417 325
rect 331 110 337 119
rect 166 52 172 90
rect 250 85 273 92
rect 250 60 257 85
rect 225 53 257 60
rect 331 59 337 102
rect 430 92 436 154
rect 495 126 501 392
rect 579 387 602 394
rect 579 362 586 387
rect 554 355 586 362
rect 660 361 666 404
rect 579 343 586 355
rect 640 354 666 361
rect 481 119 502 126
rect 395 85 436 92
rect 496 98 502 119
rect 411 60 418 85
rect 250 32 257 53
rect 311 52 357 59
rect 411 53 443 60
rect 496 57 502 90
rect 678 57 682 531
rect 250 26 303 32
rect 331 5 337 52
rect 411 29 418 53
rect 496 52 682 57
rect 994 937 1799 941
rect 994 5 999 937
rect 2068 620 2073 1666
rect 2177 1295 2183 1949
rect 2233 1929 2240 1949
rect 2300 1929 2307 1949
rect 2267 1875 2274 1891
rect 2267 1868 2318 1875
rect 2299 1843 2306 1868
rect 2233 1790 2240 1805
rect 2674 1791 2679 2445
rect 2535 1790 2563 1791
rect 2202 1784 2261 1790
rect 2269 1785 2563 1790
rect 2571 1785 2679 1791
rect 2269 1784 2542 1785
rect 2202 1460 2208 1784
rect 2233 1769 2240 1784
rect 2535 1770 2542 1784
rect 2299 1706 2306 1731
rect 2330 1706 2336 1762
rect 2601 1707 2608 1732
rect 2267 1699 2541 1706
rect 2569 1700 2632 1707
rect 2267 1683 2274 1699
rect 2233 1625 2240 1645
rect 2300 1626 2307 1645
rect 2330 1644 2336 1699
rect 2569 1684 2576 1700
rect 2535 1626 2542 1646
rect 2602 1626 2609 1646
rect 2300 1625 2425 1626
rect 2233 1619 2249 1625
rect 2257 1621 2425 1625
rect 2257 1619 2307 1621
rect 2233 1599 2240 1619
rect 2300 1599 2307 1619
rect 2356 1609 2360 1621
rect 2409 1620 2425 1621
rect 2433 1620 2551 1626
rect 2559 1620 2661 1626
rect 2267 1545 2274 1561
rect 2409 1600 2416 1620
rect 2476 1600 2483 1620
rect 2535 1600 2542 1620
rect 2602 1600 2609 1620
rect 2364 1545 2368 1559
rect 2443 1546 2450 1562
rect 2569 1546 2576 1562
rect 2629 1546 2635 1592
rect 2267 1540 2356 1545
rect 2364 1540 2417 1545
rect 2267 1538 2306 1540
rect 2299 1513 2306 1538
rect 2364 1537 2368 1540
rect 2443 1539 2543 1546
rect 2569 1539 2635 1546
rect 2356 1513 2360 1517
rect 2475 1514 2482 1539
rect 2341 1508 2390 1513
rect 2233 1460 2240 1475
rect 2341 1460 2346 1508
rect 2507 1481 2512 1539
rect 2601 1514 2608 1539
rect 2409 1461 2416 1476
rect 2535 1461 2542 1476
rect 2409 1460 2437 1461
rect 2202 1454 2261 1460
rect 2269 1455 2437 1460
rect 2445 1455 2563 1461
rect 2571 1455 2609 1461
rect 2269 1454 2410 1455
rect 2233 1439 2240 1454
rect 2299 1376 2306 1401
rect 2466 1376 2474 1405
rect 2231 1369 2474 1376
rect 2267 1353 2274 1369
rect 2233 1295 2240 1315
rect 2300 1295 2307 1315
rect 2656 1295 2661 1620
rect 2177 1289 2249 1295
rect 2257 1289 2661 1295
rect 2177 635 2183 1289
rect 2233 1269 2240 1289
rect 2300 1269 2307 1289
rect 2267 1215 2274 1231
rect 2267 1208 2318 1215
rect 2299 1183 2306 1208
rect 2233 1130 2240 1145
rect 2674 1131 2679 1785
rect 2535 1130 2563 1131
rect 2202 1124 2261 1130
rect 2269 1125 2563 1130
rect 2571 1125 2679 1131
rect 2269 1124 2542 1125
rect 2202 800 2208 1124
rect 2233 1109 2240 1124
rect 2535 1110 2542 1124
rect 2299 1046 2306 1071
rect 2330 1046 2336 1102
rect 2601 1047 2608 1072
rect 2267 1039 2541 1046
rect 2569 1040 2632 1047
rect 2267 1023 2274 1039
rect 2233 965 2240 985
rect 2300 966 2307 985
rect 2330 984 2336 1039
rect 2569 1024 2576 1040
rect 2535 966 2542 986
rect 2602 966 2609 986
rect 2300 965 2425 966
rect 2233 959 2249 965
rect 2257 961 2425 965
rect 2257 959 2307 961
rect 2233 939 2240 959
rect 2300 939 2307 959
rect 2356 949 2360 961
rect 2409 960 2425 961
rect 2433 960 2551 966
rect 2559 960 2661 966
rect 2267 885 2274 901
rect 2409 940 2416 960
rect 2476 940 2483 960
rect 2535 940 2542 960
rect 2602 940 2609 960
rect 2364 885 2368 899
rect 2443 886 2450 902
rect 2569 886 2576 902
rect 2629 886 2635 932
rect 2267 880 2356 885
rect 2364 880 2417 885
rect 2267 878 2306 880
rect 2299 853 2306 878
rect 2364 877 2368 880
rect 2443 879 2543 886
rect 2569 879 2635 886
rect 2356 853 2360 857
rect 2475 854 2482 879
rect 2341 848 2390 853
rect 2233 800 2240 815
rect 2341 800 2346 848
rect 2507 821 2512 879
rect 2601 854 2608 879
rect 2409 801 2416 816
rect 2535 801 2542 816
rect 2409 800 2437 801
rect 2202 794 2261 800
rect 2269 795 2437 800
rect 2445 795 2563 801
rect 2571 795 2609 801
rect 2269 794 2410 795
rect 2233 779 2240 794
rect 2299 716 2306 741
rect 2466 716 2474 745
rect 2231 709 2474 716
rect 2267 693 2274 709
rect 2233 635 2240 655
rect 2300 635 2307 655
rect 2656 635 2661 960
rect 2177 629 2249 635
rect 2257 629 2661 635
rect 2674 620 2679 1125
rect 2068 614 2679 620
rect 0 0 999 5
use dff_tr  dff_tr_0
timestamp 1618693583
transform 0 1 495 -1 0 3792
box -45 -495 439 171
use prop_tr1  prop_tr1_0
timestamp 1618602378
transform 1 0 697 0 1 3648
box 1 -353 386 153
<< labels >>
rlabel metal1 1064 3382 1064 3382 1 pin_p
rlabel metal1 788 3079 788 3079 1 vdd
rlabel metal1 796 3244 796 3244 5 gnd
rlabel metal1 1035 3245 1035 3245 5 gnd
rlabel metal1 1027 3080 1027 3080 1 vdd
rlabel metal1 912 3080 912 3080 1 vdd
rlabel metal1 920 3245 920 3245 5 gnd
rlabel metal1 920 2915 920 2915 1 gnd
rlabel metal1 701 2777 701 2777 3 vdd
rlabel metal1 815 2776 815 2776 7 gnd
rlabel metal1 702 2836 702 2836 3 vdd
rlabel metal1 867 2828 867 2828 7 gnd
rlabel metal1 782 2724 782 2724 1 gout2
rlabel metal1 867 2589 867 2589 7 gnd
rlabel metal1 702 2581 702 2581 3 vdd
rlabel metal1 815 2641 815 2641 7 gnd
rlabel metal1 701 2640 701 2640 3 vdd
rlabel metal1 920 2502 920 2502 5 gnd
rlabel metal1 920 2172 920 2172 1 gnd
rlabel metal1 912 2337 912 2337 5 vdd
rlabel metal1 1027 2337 1027 2337 5 vdd
rlabel metal1 1035 2172 1035 2172 1 gnd
rlabel metal1 796 2173 796 2173 1 gnd
rlabel metal1 788 2338 788 2338 5 vdd
rlabel metal1 781 2673 781 2673 1 gout3
rlabel metal1 1061 2256 1061 2256 1 pin_p3
rlabel metal1 867 1702 867 1702 7 gnd
rlabel metal1 702 1710 702 1710 3 vdd
rlabel metal1 815 1650 815 1650 7 gnd
rlabel metal1 701 1651 701 1651 3 vdd
rlabel metal1 920 1789 920 1789 1 gnd
rlabel metal1 920 2119 920 2119 5 gnd
rlabel metal1 912 1954 912 1954 1 vdd
rlabel metal1 1027 1954 1027 1954 1 vdd
rlabel metal1 1035 2119 1035 2119 5 gnd
rlabel metal1 796 2118 796 2118 5 gnd
rlabel metal1 788 1953 788 1953 1 vdd
rlabel metal1 1062 2035 1062 2035 1 pin_p4
rlabel metal1 781 1619 781 1619 1 gout4
rlabel polysilicon 793 1837 793 1837 1 A3
rlabel polysilicon 832 1938 832 1938 1 B3
rlabel polysilicon 832 2353 832 2353 1 B2
rlabel polysilicon 793 2454 793 2454 1 A2
rlabel polysilicon 793 2966 793 2966 1 A1
rlabel polysilicon 832 3059 832 3059 1 B1
rlabel metal1 333 3254 333 3254 7 vdd
rlabel metal1 3 3254 3 3254 3 vdd
rlabel metal1 168 3246 168 3246 7 gnd
rlabel metal1 169 3070 169 3070 3 gnd
rlabel metal1 334 3078 334 3078 7 vdd
rlabel polysilicon 340 3289 340 3289 3 clk
rlabel metal1 334 2952 334 2952 3 vdd
rlabel metal1 169 2956 169 2956 3 gnd
rlabel metal1 499 2950 499 2950 3 gnd
rlabel metal1 498 3246 498 3246 3 gnd
rlabel metal1 663 3254 663 3254 7 vdd
rlabel metal1 220 3176 220 3176 3 gnd
rlabel metal1 334 3177 334 3177 7 vdd
rlabel metal1 334 2698 334 2698 7 vdd
rlabel metal1 220 2697 220 2697 3 gnd
rlabel metal1 663 2775 663 2775 7 vdd
rlabel metal1 498 2767 498 2767 3 gnd
rlabel metal1 499 2471 499 2471 3 gnd
rlabel metal1 169 2477 169 2477 3 gnd
rlabel metal1 334 2473 334 2473 3 vdd
rlabel polysilicon 340 2810 340 2810 3 clk
rlabel metal1 334 2599 334 2599 7 vdd
rlabel metal1 169 2591 169 2591 3 gnd
rlabel metal1 168 2767 168 2767 7 gnd
rlabel metal1 3 2775 3 2775 3 vdd
rlabel metal1 333 2775 333 2775 7 vdd
rlabel metal1 334 2219 334 2219 7 vdd
rlabel metal1 220 2218 220 2218 3 gnd
rlabel metal1 663 2296 663 2296 7 vdd
rlabel metal1 498 2288 498 2288 3 gnd
rlabel metal1 499 1992 499 1992 3 gnd
rlabel metal1 169 1998 169 1998 3 gnd
rlabel metal1 334 1994 334 1994 3 vdd
rlabel polysilicon 340 2331 340 2331 3 clk
rlabel metal1 334 2120 334 2120 7 vdd
rlabel metal1 169 2112 169 2112 3 gnd
rlabel metal1 168 2288 168 2288 7 gnd
rlabel metal1 3 2296 3 2296 3 vdd
rlabel metal1 333 2296 333 2296 7 vdd
rlabel metal1 334 1740 334 1740 7 vdd
rlabel metal1 220 1739 220 1739 3 gnd
rlabel metal1 663 1817 663 1817 7 vdd
rlabel metal1 498 1809 498 1809 3 gnd
rlabel metal1 499 1513 499 1513 3 gnd
rlabel metal1 169 1519 169 1519 3 gnd
rlabel metal1 334 1515 334 1515 3 vdd
rlabel polysilicon 340 1852 340 1852 3 clk
rlabel metal1 334 1641 334 1641 7 vdd
rlabel metal1 169 1633 169 1633 3 gnd
rlabel metal1 168 1809 168 1809 7 gnd
rlabel metal1 3 1817 3 1817 3 vdd
rlabel metal1 333 1817 333 1817 7 vdd
rlabel metal1 333 1338 333 1338 7 vdd
rlabel metal1 3 1338 3 1338 3 vdd
rlabel metal1 168 1330 168 1330 7 gnd
rlabel metal1 169 1154 169 1154 3 gnd
rlabel metal1 334 1162 334 1162 7 vdd
rlabel polysilicon 340 1373 340 1373 3 clk
rlabel metal1 334 1036 334 1036 3 vdd
rlabel metal1 169 1040 169 1040 3 gnd
rlabel metal1 499 1034 499 1034 3 gnd
rlabel metal1 498 1330 498 1330 3 gnd
rlabel metal1 663 1338 663 1338 7 vdd
rlabel metal1 220 1260 220 1260 3 gnd
rlabel metal1 334 1261 334 1261 7 vdd
rlabel metal1 333 859 333 859 7 vdd
rlabel metal1 3 859 3 859 3 vdd
rlabel metal1 168 851 168 851 7 gnd
rlabel metal1 169 675 169 675 3 gnd
rlabel metal1 334 683 334 683 7 vdd
rlabel polysilicon 340 894 340 894 3 clk
rlabel metal1 334 557 334 557 3 vdd
rlabel metal1 169 561 169 561 3 gnd
rlabel metal1 499 555 499 555 3 gnd
rlabel metal1 498 851 498 851 3 gnd
rlabel metal1 663 859 663 859 7 vdd
rlabel metal1 220 781 220 781 3 gnd
rlabel metal1 334 782 334 782 7 vdd
rlabel metal1 333 4211 333 4211 7 vdd
rlabel metal1 3 4211 3 4211 3 vdd
rlabel metal1 168 4203 168 4203 7 gnd
rlabel metal1 169 4027 169 4027 3 gnd
rlabel metal1 334 4035 334 4035 7 vdd
rlabel polysilicon 340 4246 340 4246 3 clk
rlabel metal1 334 3909 334 3909 3 vdd
rlabel metal1 169 3913 169 3913 3 gnd
rlabel metal1 499 3907 499 3907 3 gnd
rlabel metal1 498 4203 498 4203 3 gnd
rlabel metal1 663 4211 663 4211 7 vdd
rlabel metal1 220 4133 220 4133 3 gnd
rlabel metal1 334 4134 334 4134 7 vdd
rlabel polysilicon 96 893 96 893 1 D3
rlabel polysilicon 96 1372 96 1372 1 Db2
rlabel polysilicon 96 1851 96 1851 1 D2
rlabel polysilicon 96 2330 96 2330 1 Db1
rlabel polysilicon 96 2809 96 2809 1 D1
rlabel polysilicon 179 3763 179 3763 1 clk
rlabel polysilicon 96 414 96 414 1 Db3
rlabel metal1 334 303 334 303 7 vdd
rlabel metal1 220 302 220 302 3 gnd
rlabel metal1 663 380 663 380 7 vdd
rlabel metal1 498 372 498 372 3 gnd
rlabel metal1 499 76 499 76 3 gnd
rlabel metal1 169 82 169 82 3 gnd
rlabel metal1 334 78 334 78 3 vdd
rlabel polysilicon 340 415 340 415 3 clk
rlabel metal1 334 204 334 204 7 vdd
rlabel metal1 169 196 169 196 3 gnd
rlabel metal1 168 372 168 372 7 gnd
rlabel metal1 3 380 3 380 3 vdd
rlabel metal1 333 380 333 380 7 vdd
rlabel polysilicon 96 3288 96 3288 1 carry_in
rlabel polysilicon 96 4245 96 4245 1 da0
rlabel metal1 1081 3344 1081 3344 3 gnd
rlabel metal1 1246 3352 1246 3352 7 vdd
rlabel metal1 1133 3292 1133 3292 3 gnd
rlabel metal1 1247 3293 1247 3293 7 vdd
rlabel metal1 1090 3123 1090 3123 3 gnd
rlabel metal1 1255 3131 1255 3131 7 vdd
rlabel metal1 1142 3071 1142 3071 3 gnd
rlabel metal1 1256 3072 1256 3072 7 vdd
rlabel metal1 1091 2918 1091 2918 3 gnd
rlabel metal1 1256 2926 1256 2926 7 vdd
rlabel metal1 1143 2866 1143 2866 3 gnd
rlabel metal1 1257 2867 1257 2867 7 vdd
rlabel metal1 1143 2606 1143 2606 3 gnd
rlabel metal1 1257 2605 1257 2605 7 vdd
rlabel metal1 1143 2785 1143 2785 3 gnd
rlabel metal1 1257 2786 1257 2786 7 vdd
rlabel metal1 1092 2669 1092 2669 3 gnd
rlabel metal1 1257 2677 1257 2677 7 vdd
rlabel metal1 1142 2337 1142 2337 5 vdd
rlabel metal1 1202 2224 1202 2224 1 gnd
rlabel metal1 1201 2338 1201 2338 5 vdd
rlabel metal1 1202 2120 1202 2120 5 gnd
rlabel metal1 1138 2172 1138 2172 5 gnd
rlabel metal1 1415 2556 1415 2556 7 gnd
rlabel metal1 1301 2555 1301 2555 3 vdd
rlabel metal1 1415 2735 1415 2735 7 gnd
rlabel metal1 1301 2736 1301 2736 3 vdd
rlabel metal1 1466 2619 1466 2619 7 gnd
rlabel metal1 1301 2627 1301 2627 3 vdd
rlabel metal1 1381 2599 1381 2599 1 carry_2
rlabel metal1 1142 2007 1142 2007 1 vdd
rlabel metal1 1201 2006 1201 2006 1 vdd
rlabel metal1 1201 1992 1201 1992 5 vdd
rlabel metal1 1202 1878 1202 1878 1 gnd
rlabel metal1 1142 1991 1142 1991 5 vdd
rlabel metal1 1143 1826 1143 1826 1 gnd
rlabel metal1 1478 2201 1478 2201 7 gnd
rlabel metal1 1364 2200 1364 2200 3 vdd
rlabel metal1 1478 2380 1478 2380 7 gnd
rlabel metal1 1364 2381 1364 2381 3 vdd
rlabel metal1 1529 2264 1529 2264 7 gnd
rlabel metal1 1364 2272 1364 2272 3 vdd
rlabel metal1 1482 1966 1482 1966 7 gnd
rlabel metal1 1368 1965 1368 1965 3 vdd
rlabel metal1 1482 2145 1482 2145 7 gnd
rlabel metal1 1368 2146 1368 2146 3 vdd
rlabel metal1 1533 2029 1533 2029 7 gnd
rlabel metal1 1368 2037 1368 2037 3 vdd
rlabel metal1 1594 2031 1594 2031 3 gnd
rlabel metal1 1708 2030 1708 2030 7 vdd
rlabel metal1 1594 2210 1594 2210 3 gnd
rlabel metal1 1708 2211 1708 2211 7 vdd
rlabel metal1 1543 2094 1543 2094 3 gnd
rlabel metal1 1708 2102 1708 2102 7 vdd
rlabel metal1 1628 2074 1628 2074 1 carry_3
rlabel metal1 1198 1623 1198 1623 1 vdd
rlabel metal1 1199 1737 1199 1737 5 gnd
rlabel metal1 1139 1624 1139 1624 1 vdd
rlabel metal1 1140 1789 1140 1789 5 gnd
rlabel metal1 1194 1422 1194 1422 1 vdd
rlabel metal1 1195 1536 1195 1536 5 gnd
rlabel metal1 1135 1423 1135 1423 1 vdd
rlabel metal1 1136 1588 1136 1588 5 gnd
rlabel metal1 1194 1410 1194 1410 5 vdd
rlabel metal1 1195 1296 1195 1296 1 gnd
rlabel metal1 1135 1409 1135 1409 5 vdd
rlabel metal1 1136 1244 1136 1244 1 gnd
rlabel metal1 1194 1049 1194 1049 1 vdd
rlabel metal1 1195 1163 1195 1163 5 gnd
rlabel metal1 1135 1050 1135 1050 1 vdd
rlabel metal1 1136 1215 1136 1215 5 gnd
rlabel metal1 1575 1430 1575 1430 7 gnd
rlabel metal1 1461 1429 1461 1429 3 vdd
rlabel metal1 1575 1609 1575 1609 7 gnd
rlabel metal1 1461 1610 1461 1610 3 vdd
rlabel metal1 1626 1493 1626 1493 7 gnd
rlabel metal1 1461 1501 1461 1501 3 vdd
rlabel metal1 1579 1195 1579 1195 7 gnd
rlabel metal1 1465 1194 1465 1194 3 vdd
rlabel metal1 1579 1374 1579 1374 7 gnd
rlabel metal1 1465 1375 1465 1375 3 vdd
rlabel metal1 1630 1258 1630 1258 7 gnd
rlabel metal1 1465 1266 1465 1266 3 vdd
rlabel metal1 1691 1260 1691 1260 3 gnd
rlabel metal1 1805 1259 1805 1259 7 vdd
rlabel metal1 1691 1439 1691 1439 3 gnd
rlabel metal1 1805 1440 1805 1440 7 vdd
rlabel metal1 1640 1323 1640 1323 3 gnd
rlabel metal1 1805 1331 1805 1331 7 vdd
rlabel metal1 1796 1069 1796 1069 7 vdd
rlabel metal1 1631 1061 1631 1061 3 gnd
rlabel metal1 1796 1178 1796 1178 7 vdd
rlabel metal1 1682 1177 1682 1177 3 gnd
rlabel metal1 1796 997 1796 997 7 vdd
rlabel metal1 1682 998 1682 998 3 gnd
rlabel polysilicon 1152 3343 1152 3343 1 cin0
rlabel metal1 1715 1041 1715 1041 1 carr4
rlabel metal1 1132 3446 1132 3446 3 gnd
rlabel metal1 1246 3445 1246 3445 7 vdd
rlabel metal1 1132 3625 1132 3625 3 gnd
rlabel metal1 1246 3626 1246 3626 7 vdd
rlabel metal1 1081 3509 1081 3509 3 gnd
rlabel metal1 1246 3517 1246 3517 7 vdd
rlabel metal1 2151 3336 2151 3336 3 gnd
rlabel metal1 1990 3602 1990 3602 5 gnd
rlabel metal1 1990 3272 1990 3272 1 gnd
rlabel metal1 2105 3272 2105 3272 1 gnd
rlabel metal1 2128 3356 2128 3356 1 add_out
rlabel metal1 1858 3438 1858 3438 5 vdd
rlabel metal1 2097 3437 2097 3437 5 vdd
rlabel metal1 1982 3437 1982 3437 5 vdd
rlabel metal1 1982 2960 1982 2960 1 vdd
rlabel metal1 2097 2960 2097 2960 1 vdd
rlabel metal1 1858 2959 1858 2959 1 vdd
rlabel metal1 2105 3125 2105 3125 5 gnd
rlabel metal1 1990 3125 1990 3125 5 gnd
rlabel metal1 1990 2795 1990 2795 1 gnd
rlabel metal1 2151 3061 2151 3061 3 gnd
rlabel metal1 2151 2210 2151 2210 3 gnd
rlabel metal1 1990 2476 1990 2476 5 gnd
rlabel metal1 1990 2146 1990 2146 1 gnd
rlabel metal1 2105 2146 2105 2146 1 gnd
rlabel metal1 1858 2312 1858 2312 5 vdd
rlabel metal1 2097 2311 2097 2311 5 vdd
rlabel metal1 1982 2311 1982 2311 5 vdd
rlabel metal1 2151 1935 2151 1935 3 gnd
rlabel metal1 1990 1669 1990 1669 1 gnd
rlabel metal1 1990 1999 1990 1999 5 gnd
rlabel metal1 2105 1999 2105 1999 5 gnd
rlabel metal1 1858 1833 1858 1833 1 vdd
rlabel metal1 2097 1834 2097 1834 1 vdd
rlabel metal1 1982 1834 1982 1834 1 vdd
rlabel polysilicon 1871 3189 1871 3189 1 cin1
rlabel polysilicon 1871 2082 1871 2082 1 cin2
rlabel metal1 2128 1915 2128 1915 1 add_out3
rlabel metal1 2128 2230 2128 2230 1 add_out2
rlabel metal1 2128 3041 2128 3041 1 add_out1
rlabel metal1 2281 2942 2281 2942 5 vdd
rlabel metal1 2289 2777 2289 2777 5 gnd
rlabel metal1 2465 2778 2465 2778 1 gnd
rlabel metal1 2457 2943 2457 2943 5 vdd
rlabel polysilicon 2246 2949 2246 2949 1 clk
rlabel metal1 2583 2943 2583 2943 1 vdd
rlabel metal1 2579 2778 2579 2778 1 gnd
rlabel metal1 2585 3108 2585 3108 1 gnd
rlabel metal1 2289 3107 2289 3107 1 gnd
rlabel metal1 2359 2829 2359 2829 1 gnd
rlabel metal1 2358 2943 2358 2943 5 vdd
rlabel metal1 2281 2282 2281 2282 5 vdd
rlabel metal1 2289 2117 2289 2117 5 gnd
rlabel metal1 2465 2118 2465 2118 1 gnd
rlabel metal1 2457 2283 2457 2283 5 vdd
rlabel polysilicon 2246 2289 2246 2289 1 clk
rlabel metal1 2583 2283 2583 2283 1 vdd
rlabel metal1 2579 2118 2579 2118 1 gnd
rlabel metal1 2585 2448 2585 2448 1 gnd
rlabel metal1 2289 2447 2289 2447 1 gnd
rlabel metal1 2281 2612 2281 2612 5 vdd
rlabel metal1 2359 2169 2359 2169 1 gnd
rlabel metal1 2358 2283 2358 2283 5 vdd
rlabel metal1 2281 1622 2281 1622 5 vdd
rlabel metal1 2289 1457 2289 1457 5 gnd
rlabel metal1 2465 1458 2465 1458 1 gnd
rlabel metal1 2457 1623 2457 1623 5 vdd
rlabel polysilicon 2246 1629 2246 1629 1 clk
rlabel metal1 2583 1623 2583 1623 1 vdd
rlabel metal1 2579 1458 2579 1458 1 gnd
rlabel metal1 2585 1788 2585 1788 1 gnd
rlabel metal1 2289 1787 2289 1787 1 gnd
rlabel metal1 2281 1952 2281 1952 5 vdd
rlabel metal1 2359 1509 2359 1509 1 gnd
rlabel metal1 2358 1623 2358 1623 5 vdd
rlabel metal1 2281 962 2281 962 5 vdd
rlabel metal1 2289 797 2289 797 5 gnd
rlabel metal1 2465 798 2465 798 1 gnd
rlabel metal1 2457 963 2457 963 5 vdd
rlabel polysilicon 2246 969 2246 969 1 clk
rlabel metal1 2583 963 2583 963 1 vdd
rlabel metal1 2579 798 2579 798 1 gnd
rlabel metal1 2585 1128 2585 1128 1 gnd
rlabel metal1 2289 1127 2289 1127 1 gnd
rlabel metal1 2281 1292 2281 1292 5 vdd
rlabel metal1 2359 849 2359 849 1 gnd
rlabel metal1 2358 963 2358 963 5 vdd
rlabel metal1 2281 632 2281 632 5 vdd
rlabel metal1 2627 3023 2627 3023 1 sum_1
rlabel metal1 2631 2862 2631 2862 1 sum_1_bar
rlabel metal1 2627 2363 2627 2363 1 sum_2
rlabel metal1 2631 2202 2631 2202 1 sum_2_bar
rlabel metal1 2627 1703 2627 1703 1 sum_3
rlabel metal1 2630 1542 2630 1542 1 sum_3_bar
rlabel metal1 2627 1043 2627 1043 1 carry_4
rlabel metal1 2631 882 2631 882 1 carry_4_bar
rlabel metal1 2358 3603 2358 3603 5 vdd
rlabel metal1 2359 3489 2359 3489 1 gnd
rlabel metal1 2281 3932 2281 3932 5 vdd
rlabel metal1 2289 3767 2289 3767 1 gnd
rlabel metal1 2585 3768 2585 3768 1 gnd
rlabel metal1 2579 3438 2579 3438 1 gnd
rlabel metal1 2583 3603 2583 3603 1 vdd
rlabel metal1 2457 3603 2457 3603 5 vdd
rlabel metal1 2465 3438 2465 3438 1 gnd
rlabel metal1 2289 3437 2289 3437 5 gnd
rlabel metal1 2281 3272 2281 3272 1 vdd
rlabel metal1 2281 3602 2281 3602 5 vdd
rlabel metal1 2630 3523 2630 3523 1 sum_0_bar
rlabel metal1 2629 3684 2629 3684 1 sum_out
rlabel metal1 2510 3522 2510 3522 1 dfo1
rlabel metal1 2338 3353 2338 3353 1 dfo2
rlabel polysilicon 2550 3682 2550 3682 1 dfi1
rlabel polysilicon 2592 3697 2592 3697 1 dfi2
rlabel polysilicon 2553 3507 2553 3507 1 din3
rlabel polysilicon 2246 3610 2246 3610 1 clk
<< end >>
