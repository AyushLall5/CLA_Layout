magic
tech scmos
timestamp 1618606384
<< nwell >>
rect 699 227 796 283
rect 575 148 672 204
rect 699 147 796 203
rect 814 147 911 203
rect 473 109 552 134
rect 480 0 536 97
<< ntransistor >>
rect 727 324 729 364
rect 766 324 768 364
rect 443 121 463 123
rect 399 67 439 69
rect 603 67 605 107
rect 642 67 644 107
rect 399 28 439 30
rect 727 66 729 106
rect 766 66 768 106
rect 842 66 844 106
rect 881 66 883 106
<< ptransistor >>
rect 727 236 729 276
rect 766 236 768 276
rect 603 155 605 195
rect 642 155 644 195
rect 485 121 535 123
rect 727 154 729 194
rect 766 154 768 194
rect 842 154 844 194
rect 881 154 883 194
rect 487 67 527 69
rect 487 28 527 30
<< ndiffusion >>
rect 707 362 727 364
rect 707 324 710 362
rect 717 324 727 362
rect 729 324 766 364
rect 768 362 787 364
rect 768 324 776 362
rect 783 324 787 362
rect 443 123 463 124
rect 443 120 463 121
rect 399 84 439 88
rect 399 77 401 84
rect 399 69 439 77
rect 583 69 586 107
rect 593 69 603 107
rect 583 67 603 69
rect 605 67 642 107
rect 644 69 652 107
rect 659 69 663 107
rect 644 67 663 69
rect 707 68 710 106
rect 717 68 727 106
rect 399 30 439 67
rect 399 18 439 28
rect 399 11 401 18
rect 399 8 439 11
rect 707 66 727 68
rect 729 66 766 106
rect 768 68 776 106
rect 783 68 787 106
rect 768 66 787 68
rect 822 68 825 106
rect 832 68 842 106
rect 822 66 842 68
rect 844 66 881 106
rect 883 68 891 106
rect 898 68 902 106
rect 883 66 902 68
<< pdiffusion >>
rect 707 238 710 276
rect 717 238 727 276
rect 707 236 727 238
rect 729 238 744 276
rect 751 238 766 276
rect 729 236 766 238
rect 768 238 777 276
rect 784 238 787 276
rect 768 236 787 238
rect 583 193 603 195
rect 583 155 586 193
rect 593 155 603 193
rect 605 193 642 195
rect 605 155 620 193
rect 627 155 642 193
rect 644 193 663 195
rect 644 155 653 193
rect 660 155 663 193
rect 485 123 535 124
rect 485 120 535 121
rect 707 192 727 194
rect 707 154 710 192
rect 717 154 727 192
rect 729 192 766 194
rect 729 154 744 192
rect 751 154 766 192
rect 768 192 787 194
rect 768 154 777 192
rect 784 154 787 192
rect 822 192 842 194
rect 822 154 825 192
rect 832 154 842 192
rect 844 192 881 194
rect 844 154 859 192
rect 866 154 881 192
rect 883 192 902 194
rect 883 154 892 192
rect 899 154 902 192
rect 487 85 527 88
rect 525 78 527 85
rect 487 69 527 78
rect 487 52 527 67
rect 525 45 527 52
rect 487 30 527 45
rect 487 18 527 28
rect 525 11 527 18
rect 487 8 527 11
<< ndcontact >>
rect 710 324 717 362
rect 776 324 783 362
rect 443 124 463 128
rect 443 116 463 120
rect 401 77 439 84
rect 586 69 593 107
rect 652 69 659 107
rect 710 68 717 106
rect 401 11 439 18
rect 776 68 783 106
rect 825 68 832 106
rect 891 68 898 106
<< pdcontact >>
rect 710 238 717 276
rect 744 238 751 276
rect 777 238 784 276
rect 586 155 593 193
rect 620 155 627 193
rect 653 155 660 193
rect 485 124 535 128
rect 485 116 535 120
rect 710 154 717 192
rect 744 154 751 192
rect 777 154 784 192
rect 825 154 832 192
rect 859 154 866 192
rect 892 154 899 192
rect 487 78 525 85
rect 487 45 525 52
rect 487 11 525 18
<< psubstratepcontact >>
rect 738 377 746 383
rect 380 39 386 47
rect 614 48 622 54
rect 738 47 746 53
rect 853 47 861 53
<< nsubstratencontact >>
rect 602 213 610 219
rect 726 212 734 218
rect 841 212 849 218
rect 545 27 551 35
<< polysilicon >>
rect 727 364 729 367
rect 766 364 768 367
rect 727 294 729 324
rect 623 292 729 294
rect 623 209 625 292
rect 727 276 729 292
rect 766 276 768 324
rect 876 294 883 296
rect 727 233 729 236
rect 766 225 768 236
rect 603 207 625 209
rect 686 223 768 225
rect 603 195 605 207
rect 642 195 644 198
rect 440 121 443 123
rect 463 121 485 123
rect 535 121 538 123
rect 603 107 605 155
rect 642 117 644 155
rect 686 139 688 223
rect 727 194 729 197
rect 766 194 768 197
rect 842 194 844 197
rect 881 194 883 294
rect 727 117 729 154
rect 766 126 768 154
rect 842 135 844 154
rect 834 133 844 135
rect 760 124 768 126
rect 642 115 729 117
rect 642 107 644 115
rect 373 86 392 88
rect 390 69 392 86
rect 390 67 399 69
rect 439 67 487 69
rect 527 67 542 69
rect 727 106 729 115
rect 766 106 768 124
rect 842 106 844 133
rect 881 106 883 154
rect 540 63 542 67
rect 603 63 605 67
rect 540 61 605 63
rect 396 28 399 30
rect 439 28 487 30
rect 527 28 530 30
rect 456 -13 458 28
rect 642 -13 644 67
rect 727 63 729 66
rect 766 63 768 66
rect 842 63 844 66
rect 881 63 883 66
rect 456 -15 644 -13
<< polycontact >>
rect 871 292 876 299
rect 466 116 471 121
rect 684 134 691 139
rect 756 122 760 128
rect 829 131 834 138
rect 368 83 373 91
<< metal1 >>
rect 0 537 562 542
rect 0 486 5 537
rect 81 521 481 527
rect 81 500 86 521
rect 476 375 481 521
rect 557 365 562 537
rect 710 377 738 383
rect 746 377 929 383
rect 710 362 717 377
rect 776 299 783 324
rect 744 292 871 299
rect 744 276 751 292
rect 484 261 489 262
rect 710 219 717 238
rect 475 215 482 219
rect 561 213 602 219
rect 610 218 717 219
rect 777 218 784 238
rect 610 213 726 218
rect 384 178 392 205
rect 586 193 593 213
rect 653 212 726 213
rect 734 212 841 218
rect 849 212 899 218
rect 653 193 660 212
rect 476 156 481 161
rect 466 152 481 156
rect 434 120 439 150
rect 466 128 471 152
rect 557 134 562 168
rect 710 192 717 212
rect 777 192 784 212
rect 547 129 562 134
rect 620 139 627 155
rect 825 192 832 212
rect 892 192 899 212
rect 620 132 659 139
rect 463 124 485 128
rect 434 116 443 120
rect 547 120 552 129
rect 535 116 552 120
rect 434 106 439 116
rect 380 101 439 106
rect 361 83 368 91
rect 380 47 386 101
rect 466 84 471 116
rect 547 85 552 116
rect 652 128 659 132
rect 684 128 691 134
rect 744 138 751 154
rect 859 138 866 154
rect 744 131 829 138
rect 859 131 907 138
rect 652 122 756 128
rect 652 107 659 122
rect 439 77 471 84
rect 525 78 552 85
rect 464 52 471 77
rect 464 45 487 52
rect 380 18 386 39
rect 545 35 552 78
rect 776 106 783 131
rect 891 106 898 131
rect 586 54 593 69
rect 710 54 717 68
rect 586 48 614 54
rect 622 53 717 54
rect 825 53 832 68
rect 924 53 929 377
rect 622 48 738 53
rect 551 27 552 35
rect 545 18 552 27
rect 380 11 401 18
rect 525 11 552 18
rect 380 -21 386 11
rect 545 0 552 11
rect 677 -21 683 48
rect 710 47 738 48
rect 746 47 853 53
rect 861 47 929 53
rect 380 -26 683 -21
use prop_tr1  prop_tr1_0
timestamp 1618602378
transform 1 0 -1 0 1 353
box 1 -353 386 153
use or_tr2  or_tr2_0
timestamp 1618345886
transform 0 1 391 -1 0 307
box -70 0 147 171
<< labels >>
rlabel metal1 383 67 383 67 3 gnd
rlabel metal1 435 119 435 119 3 gnd
rlabel metal1 468 148 468 148 1 o_ca
rlabel metal1 366 87 366 87 1 pin_p
rlabel metal1 478 216 478 216 1 carr_out
rlabel metal1 927 114 927 114 3 gnd
rlabel metal1 766 380 766 380 5 gnd
rlabel metal1 766 50 766 50 1 gnd
rlabel metal1 881 50 881 50 1 gnd
rlabel polysilicon 567 -14 567 -14 1 cin0
rlabel metal1 904 134 904 134 1 add_out
rlabel metal1 549 118 549 118 7 vdd
rlabel metal1 548 59 548 59 7 vdd
rlabel metal1 634 216 634 216 5 vdd
rlabel metal1 873 215 873 215 5 vdd
rlabel metal1 758 215 758 215 5 vdd
<< end >>
