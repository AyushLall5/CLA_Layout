magic
tech scmos
timestamp 1618693583
<< nwell >>
rect 0 -150 97 -94
rect 302 -149 399 -93
rect 0 -230 97 -174
rect 176 -229 273 -173
rect 302 -229 399 -173
rect 0 -480 97 -424
<< ntransistor >>
rect 28 -53 30 -13
rect 67 -53 69 -13
rect 330 -52 332 -12
rect 369 -52 371 -12
rect 28 -311 30 -271
rect 67 -311 69 -271
rect 204 -310 206 -270
rect 243 -310 245 -270
rect 28 -383 30 -343
rect 67 -383 69 -343
rect 330 -310 332 -270
rect 369 -310 371 -270
<< ptransistor >>
rect 28 -141 30 -101
rect 67 -141 69 -101
rect 330 -140 332 -100
rect 369 -140 371 -100
rect 28 -223 30 -183
rect 67 -223 69 -183
rect 204 -222 206 -182
rect 243 -222 245 -182
rect 330 -222 332 -182
rect 369 -222 371 -182
rect 28 -471 30 -431
rect 67 -471 69 -431
<< ndiffusion >>
rect 8 -15 28 -13
rect 8 -53 11 -15
rect 18 -53 28 -15
rect 30 -53 67 -13
rect 69 -15 88 -13
rect 69 -53 77 -15
rect 84 -53 88 -15
rect 310 -14 330 -12
rect 310 -52 313 -14
rect 320 -52 330 -14
rect 332 -52 369 -12
rect 371 -14 390 -12
rect 371 -52 379 -14
rect 386 -52 390 -14
rect 8 -309 11 -271
rect 18 -309 28 -271
rect 8 -311 28 -309
rect 30 -311 67 -271
rect 69 -309 77 -271
rect 84 -309 88 -271
rect 69 -311 88 -309
rect 184 -308 187 -270
rect 194 -308 204 -270
rect 184 -310 204 -308
rect 206 -310 243 -270
rect 245 -308 253 -270
rect 260 -308 264 -270
rect 245 -310 264 -308
rect 8 -345 28 -343
rect 8 -383 11 -345
rect 18 -383 28 -345
rect 30 -383 67 -343
rect 69 -345 88 -343
rect 69 -383 77 -345
rect 84 -383 88 -345
rect 310 -308 313 -270
rect 320 -308 330 -270
rect 310 -310 330 -308
rect 332 -310 369 -270
rect 371 -308 379 -270
rect 386 -308 390 -270
rect 371 -310 390 -308
<< pdiffusion >>
rect 8 -139 11 -101
rect 18 -139 28 -101
rect 8 -141 28 -139
rect 30 -139 45 -101
rect 52 -139 67 -101
rect 30 -141 67 -139
rect 69 -139 78 -101
rect 85 -139 88 -101
rect 69 -141 88 -139
rect 310 -138 313 -100
rect 320 -138 330 -100
rect 310 -140 330 -138
rect 332 -138 347 -100
rect 354 -138 369 -100
rect 332 -140 369 -138
rect 371 -138 380 -100
rect 387 -138 390 -100
rect 371 -140 390 -138
rect 8 -185 28 -183
rect 8 -223 11 -185
rect 18 -223 28 -185
rect 30 -185 67 -183
rect 30 -223 45 -185
rect 52 -223 67 -185
rect 69 -185 88 -183
rect 69 -223 78 -185
rect 85 -223 88 -185
rect 184 -184 204 -182
rect 184 -222 187 -184
rect 194 -222 204 -184
rect 206 -184 243 -182
rect 206 -222 221 -184
rect 228 -222 243 -184
rect 245 -184 264 -182
rect 245 -222 254 -184
rect 261 -222 264 -184
rect 310 -184 330 -182
rect 310 -222 313 -184
rect 320 -222 330 -184
rect 332 -184 369 -182
rect 332 -222 347 -184
rect 354 -222 369 -184
rect 371 -184 390 -182
rect 371 -222 380 -184
rect 387 -222 390 -184
rect 8 -469 11 -431
rect 18 -469 28 -431
rect 8 -471 28 -469
rect 30 -469 45 -431
rect 52 -469 67 -431
rect 30 -471 67 -469
rect 69 -469 78 -431
rect 85 -469 88 -431
rect 69 -471 88 -469
<< ndcontact >>
rect 11 -53 18 -15
rect 77 -53 84 -15
rect 313 -52 320 -14
rect 379 -52 386 -14
rect 11 -309 18 -271
rect 77 -309 84 -271
rect 187 -308 194 -270
rect 253 -308 260 -270
rect 11 -383 18 -345
rect 77 -383 84 -345
rect 313 -308 320 -270
rect 379 -308 386 -270
<< pdcontact >>
rect 11 -139 18 -101
rect 45 -139 52 -101
rect 78 -139 85 -101
rect 313 -138 320 -100
rect 347 -138 354 -100
rect 380 -138 387 -100
rect 11 -223 18 -185
rect 45 -223 52 -185
rect 78 -223 85 -185
rect 187 -222 194 -184
rect 221 -222 228 -184
rect 254 -222 261 -184
rect 313 -222 320 -184
rect 347 -222 354 -184
rect 380 -222 387 -184
rect 11 -469 18 -431
rect 45 -469 52 -431
rect 78 -469 85 -431
<< psubstratepcontact >>
rect 39 0 47 6
rect 341 1 349 7
rect 39 -330 47 -324
rect 215 -329 223 -323
rect 341 -329 349 -323
<< nsubstratencontact >>
rect 27 -165 35 -159
rect 203 -164 211 -158
rect 329 -164 337 -158
rect 27 -495 35 -489
<< polysilicon >>
rect 69 95 112 97
rect -7 80 28 82
rect -7 -410 -5 80
rect 98 -5 100 84
rect 67 -7 100 -5
rect 28 -13 30 -10
rect 67 -13 69 -7
rect 110 -17 112 95
rect 330 -12 332 -9
rect 369 -12 371 -9
rect 28 -101 30 -53
rect 67 -101 69 -53
rect 330 -81 332 -52
rect 324 -83 332 -81
rect 330 -100 332 -83
rect 369 -100 371 -52
rect 415 -81 422 -79
rect 28 -153 30 -141
rect 67 -144 69 -141
rect 330 -143 332 -140
rect 23 -155 30 -153
rect 23 -168 25 -155
rect 23 -170 30 -168
rect 110 -169 112 -147
rect 369 -152 371 -140
rect 369 -154 411 -152
rect 28 -183 30 -170
rect 67 -171 112 -169
rect 67 -183 69 -171
rect 204 -182 206 -179
rect 243 -182 245 -179
rect 330 -182 332 -179
rect 369 -182 371 -179
rect 409 -187 411 -154
rect 28 -271 30 -223
rect 67 -271 69 -223
rect 204 -240 206 -222
rect 199 -242 206 -240
rect 204 -270 206 -242
rect 243 -270 245 -222
rect 330 -241 332 -222
rect 326 -243 332 -241
rect 330 -270 332 -243
rect 369 -256 371 -222
rect 420 -256 422 -81
rect 369 -258 422 -256
rect 369 -270 371 -258
rect 28 -314 30 -311
rect 67 -314 69 -311
rect 204 -313 206 -310
rect 243 -318 245 -310
rect 243 -320 248 -318
rect 28 -343 30 -340
rect 67 -343 69 -340
rect 246 -373 248 -320
rect 28 -398 30 -383
rect 24 -400 30 -398
rect -7 -412 3 -410
rect 28 -431 30 -400
rect 67 -393 69 -383
rect 286 -393 288 -307
rect 330 -313 332 -310
rect 369 -313 371 -310
rect 67 -395 288 -393
rect 67 -431 69 -395
rect 28 -474 30 -471
rect 67 -474 69 -471
<< polycontact >>
rect 96 84 103 91
rect 108 -22 114 -17
rect 319 -85 324 -78
rect 410 -84 415 -77
rect 108 -147 114 -140
rect 407 -192 413 -187
rect 195 -244 199 -239
rect 321 -245 326 -238
rect 285 -307 290 -303
rect 244 -379 252 -373
rect 3 -415 9 -408
<< metal1 >>
rect -45 165 11 171
rect -45 -489 -39 165
rect 83 84 96 91
rect 313 6 341 7
rect -20 0 39 6
rect 47 1 341 6
rect 349 1 387 7
rect 47 0 320 1
rect -20 -324 -14 0
rect 11 -15 18 0
rect 313 -14 320 0
rect 77 -78 84 -53
rect 108 -78 114 -22
rect 379 -77 386 -52
rect 45 -85 319 -78
rect 347 -84 410 -77
rect 45 -101 52 -85
rect 11 -159 18 -139
rect 78 -158 85 -139
rect 108 -140 114 -85
rect 347 -100 354 -84
rect 313 -158 320 -138
rect 380 -158 387 -138
rect 78 -159 127 -158
rect 11 -165 27 -159
rect 35 -163 127 -159
rect 152 -163 203 -158
rect 35 -165 85 -163
rect 11 -185 18 -165
rect 78 -185 85 -165
rect 187 -164 203 -163
rect 211 -164 329 -158
rect 337 -164 439 -158
rect 187 -184 194 -164
rect 254 -184 261 -164
rect 313 -184 320 -164
rect 380 -184 387 -164
rect 45 -239 52 -223
rect 221 -238 228 -222
rect 347 -238 354 -222
rect 407 -238 413 -192
rect 45 -244 120 -239
rect 168 -244 195 -239
rect 45 -246 84 -244
rect 221 -245 321 -238
rect 347 -245 413 -238
rect 77 -271 84 -246
rect 253 -270 260 -245
rect 11 -324 18 -309
rect 119 -324 124 -276
rect 285 -303 290 -245
rect 379 -270 386 -245
rect 187 -323 194 -308
rect 313 -323 320 -308
rect 187 -324 215 -323
rect -20 -330 39 -324
rect 47 -329 215 -324
rect 223 -329 341 -323
rect 349 -329 387 -323
rect 47 -330 188 -329
rect 11 -345 18 -330
rect 77 -408 84 -383
rect 244 -408 252 -379
rect 9 -415 252 -408
rect 45 -431 52 -415
rect 11 -489 18 -469
rect 78 -489 85 -469
rect 434 -489 439 -164
rect -45 -495 27 -489
rect 35 -495 439 -489
use nand_tr  nand_tr_0
timestamp 1618160895
transform 1 0 0 0 1 100
box 0 -100 97 71
use first  first_0
timestamp 1618336112
transform 1 0 41 0 1 -233
box 78 -43 127 75
<< labels >>
rlabel metal1 67 3 67 3 5 gnd
rlabel metal1 59 -162 59 -162 5 vdd
rlabel metal1 59 -492 59 -492 1 vdd
rlabel metal1 67 -327 67 -327 5 gnd
rlabel metal1 243 -326 243 -326 1 gnd
rlabel metal1 235 -161 235 -161 5 vdd
rlabel polysilicon 24 -155 24 -155 1 clk
rlabel polysilicon 25 -399 25 -399 1 D
rlabel metal1 361 -161 361 -161 1 vdd
rlabel metal1 410 -241 410 -241 7 S_bar
rlabel metal1 357 -326 357 -326 1 gnd
rlabel metal1 405 -81 405 -81 1 S
rlabel metal1 363 4 363 4 1 gnd
<< end >>
