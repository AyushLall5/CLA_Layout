magic
tech scmos
timestamp 1618160895
<< nwell >>
rect 0 0 97 56
<< ntransistor >>
rect 28 -81 30 -41
rect 67 -81 69 -41
<< ptransistor >>
rect 28 7 30 47
rect 67 7 69 47
<< ndiffusion >>
rect 8 -79 11 -41
rect 18 -79 28 -41
rect 8 -81 28 -79
rect 30 -81 67 -41
rect 69 -79 77 -41
rect 84 -79 88 -41
rect 69 -81 88 -79
<< pdiffusion >>
rect 8 45 28 47
rect 8 7 11 45
rect 18 7 28 45
rect 30 45 67 47
rect 30 7 45 45
rect 52 7 67 45
rect 69 45 88 47
rect 69 7 78 45
rect 85 7 88 45
<< ndcontact >>
rect 11 -79 18 -41
rect 77 -79 84 -41
<< pdcontact >>
rect 11 7 18 45
rect 45 7 52 45
rect 78 7 85 45
<< psubstratepcontact >>
rect 39 -100 47 -94
<< nsubstratencontact >>
rect 27 65 35 71
<< polysilicon >>
rect 28 47 30 50
rect 67 47 69 50
rect 28 -41 30 7
rect 67 -41 69 7
rect 28 -84 30 -81
rect 67 -84 69 -81
<< metal1 >>
rect 11 65 27 71
rect 35 65 85 71
rect 11 45 18 65
rect 78 45 85 65
rect 45 -9 52 7
rect 45 -16 84 -9
rect 77 -41 84 -16
rect 11 -94 18 -79
rect 11 -100 39 -94
rect 47 -100 85 -94
<< labels >>
rlabel metal1 67 -97 67 -97 1 gnd
rlabel metal1 59 68 59 68 5 vdd
<< end >>
